// system.v

// Generated using ACDS version 14.0 200 at 2021.03.08.12:40:36

`timescale 1 ps / 1 ps
module system (
		input  wire        clk_sys_clk,                    //             clk_sys.clk
		input  wire        reset_sys_reset_n,              //           reset_sys.reset_n
		input  wire        clk_vga_clk,                    //             clk_vga.clk
		input  wire        reset_vga_reset_n,              //           reset_vga.reset_n
		output wire [12:0] sdram_conduit_end_addr,         //   sdram_conduit_end.addr
		output wire [1:0]  sdram_conduit_end_ba,           //                    .ba
		output wire        sdram_conduit_end_cas_n,        //                    .cas_n
		output wire        sdram_conduit_end_cke,          //                    .cke
		output wire        sdram_conduit_end_cs_n,         //                    .cs_n
		inout  wire [31:0] sdram_conduit_end_dq,           //                    .dq
		output wire [3:0]  sdram_conduit_end_dqm,          //                    .dqm
		output wire        sdram_conduit_end_ras_n,        //                    .ras_n
		output wire        sdram_conduit_end_we_n,         //                    .we_n
		input  wire        clk_sound_clk,                  //           clk_sound.clk
		input  wire        reset_sound_reset_n,            //         reset_sound.reset_n
		input  wire [7:0]  pio_input_export,               //           pio_input.export
		input  wire        reset_only_ao486_reset,         //    reset_only_ao486.reset
		output wire [7:0]  pio_output_export,              //          pio_output.export
		output wire        export_sound_sclk,              //        export_sound.sclk
		inout  wire        export_sound_sdat,              //                    .sdat
		output wire        export_sound_xclk,              //                    .xclk
		output wire        export_sound_bclk,              //                    .bclk
		output wire        export_sound_dat,               //                    .dat
		output wire        export_sound_lr,                //                    .lr
		output wire        export_vga_clock,               //          export_vga.clock
		output wire        export_vga_sync_n,              //                    .sync_n
		output wire        export_vga_blank_n,             //                    .blank_n
		output wire        export_vga_horiz_sync,          //                    .horiz_sync
		output wire        export_vga_vert_sync,           //                    .vert_sync
		output wire [7:0]  export_vga_r,                   //                    .r
		output wire [7:0]  export_vga_g,                   //                    .g
		output wire [7:0]  export_vga_b,                   //                    .b
		inout  wire        export_ps2_kbclk,               //          export_ps2.kbclk
		inout  wire        export_ps2_kbdat,               //                    .kbdat
		inout  wire        export_ps2_mouseclk,            //                    .mouseclk
		inout  wire        export_ps2_mousedat,            //                    .mousedat
		output wire        export_ps2_out_port_a20_enable, // export_ps2_out_port.a20_enable
		output wire        export_ps2_out_port_reset_n,    //                    .reset_n
		inout  wire [3:0]  sd_dat_export,                  //              sd_dat.export
		inout  wire        sd_cmd_export,                  //              sd_cmd.export
		output wire        sd_clk_export                   //              sd_clk.export
	);

	wire   [7:0] floppy_conduit_ide_3f6_writedata;                          // floppy:ide_3f6_writedata -> hdd:ide_3f6_writedata
	wire         floppy_conduit_ide_3f6_write;                              // floppy:ide_3f6_write -> hdd:ide_3f6_write
	wire         floppy_conduit_ide_3f6_read;                               // floppy:ide_3f6_read -> hdd:ide_3f6_read
	wire   [7:0] hdd_conduit_ide_3f6_readdata;                              // hdd:ide_3f6_readdata -> floppy:ide_3f6_readdata
	wire         pc_dma_conduit_dma_floppy_terminal;                        // pc_dma:dma_floppy_terminal -> floppy:dma_floppy_terminal
	wire   [7:0] floppy_conduit_dma_floppy_writedata;                       // floppy:dma_floppy_writedata -> pc_dma:dma_floppy_writedata
	wire         pc_dma_conduit_dma_floppy_ack;                             // pc_dma:dma_floppy_ack -> floppy:dma_floppy_ack
	wire   [7:0] pc_dma_conduit_dma_floppy_readdata;                        // pc_dma:dma_floppy_readdata -> floppy:dma_floppy_readdata
	wire         floppy_conduit_dma_floppy_req;                             // floppy:dma_floppy_req -> pc_dma:dma_floppy_req
	wire         pc_dma_conduit_dma_soundblaster_terminal;                  // pc_dma:dma_soundblaster_terminal -> sound:dma_soundblaster_terminal
	wire   [7:0] sound_conduit_dma_soundblaster_writedata;                  // sound:dma_soundblaster_writedata -> pc_dma:dma_soundblaster_writedata
	wire         pc_dma_conduit_dma_soundblaster_ack;                       // pc_dma:dma_soundblaster_ack -> sound:dma_soundblaster_ack
	wire   [7:0] pc_dma_conduit_dma_soundblaster_readdata;                  // pc_dma:dma_soundblaster_readdata -> sound:dma_soundblaster_readdata
	wire         sound_conduit_dma_soundblaster_req;                        // sound:dma_soundblaster_req -> pc_dma:dma_soundblaster_req
	wire         nios2_jtag_debug_module_reset_reset;                       // nios2:jtag_debug_module_resetrequest -> reset_sys:reset_in1
	wire         reset_sys_reset_out_reset;                                 // reset_sys:reset_out -> [reset_only_ao486:reset_in1, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	wire         pic_conduit_interrupt_interrupt_do;                        // pic:interrupt_do -> ao486:interrupt_do
	wire   [7:0] pic_conduit_interrupt_interrupt_vector;                    // pic:interrupt_vector -> ao486:interrupt_vector
	wire         ao486_interrupt_interrupt_done;                            // ao486:interrupt_done -> pic:interrupt_done
	wire         pit_conduit_speaker_enable;                                // pit:speaker_enable -> sound:speaker_enable
	wire         pit_conduit_speaker_out;                                   // pit:speaker_out -> sound:speaker_out
	wire   [7:0] ps2_conduit_speaker_61h_writedata;                         // ps2:speaker_61h_writedata -> pit:speaker_61h_writedata
	wire         ps2_conduit_speaker_61h_write;                             // ps2:speaker_61h_write -> pit:speaker_61h_write
	wire         ps2_conduit_speaker_61h_read;                              // ps2:speaker_61h_read -> pit:speaker_61h_read
	wire   [7:0] pit_conduit_speaker_61h_readdata;                          // pit:speaker_61h_readdata -> ps2:speaker_61h_readdata
	wire         reset_only_ao486_reset_out_reset;                          // reset_only_ao486:reset_out -> [ao486:rst_n, mm_interconnect_0:ao486_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:ao486_reset_sink_reset_bridge_in_reset_reset]
	wire         nios2_data_master_waitrequest;                             // mm_interconnect_0:nios2_data_master_waitrequest -> nios2:d_waitrequest
	wire  [31:0] nios2_data_master_writedata;                               // nios2:d_writedata -> mm_interconnect_0:nios2_data_master_writedata
	wire  [27:0] nios2_data_master_address;                                 // nios2:d_address -> mm_interconnect_0:nios2_data_master_address
	wire         nios2_data_master_write;                                   // nios2:d_write -> mm_interconnect_0:nios2_data_master_write
	wire         nios2_data_master_read;                                    // nios2:d_read -> mm_interconnect_0:nios2_data_master_read
	wire  [31:0] nios2_data_master_readdata;                                // mm_interconnect_0:nios2_data_master_readdata -> nios2:d_readdata
	wire         nios2_data_master_debugaccess;                             // nios2:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:nios2_data_master_debugaccess
	wire   [3:0] nios2_data_master_byteenable;                              // nios2:d_byteenable -> mm_interconnect_0:nios2_data_master_byteenable
	wire         floppy_avalon_master_waitrequest;                          // mm_interconnect_0:floppy_avalon_master_waitrequest -> floppy:sd_master_waitrequest
	wire  [31:0] floppy_avalon_master_writedata;                            // floppy:sd_master_writedata -> mm_interconnect_0:floppy_avalon_master_writedata
	wire  [31:0] floppy_avalon_master_address;                              // floppy:sd_master_address -> mm_interconnect_0:floppy_avalon_master_address
	wire         floppy_avalon_master_write;                                // floppy:sd_master_write -> mm_interconnect_0:floppy_avalon_master_write
	wire         floppy_avalon_master_read;                                 // floppy:sd_master_read -> mm_interconnect_0:floppy_avalon_master_read
	wire  [31:0] floppy_avalon_master_readdata;                             // mm_interconnect_0:floppy_avalon_master_readdata -> floppy:sd_master_readdata
	wire         floppy_avalon_master_readdatavalid;                        // mm_interconnect_0:floppy_avalon_master_readdatavalid -> floppy:sd_master_readdatavalid
	wire         hdd_avalon_master_waitrequest;                             // mm_interconnect_0:hdd_avalon_master_waitrequest -> hdd:sd_master_waitrequest
	wire  [31:0] hdd_avalon_master_writedata;                               // hdd:sd_master_writedata -> mm_interconnect_0:hdd_avalon_master_writedata
	wire  [31:0] hdd_avalon_master_address;                                 // hdd:sd_master_address -> mm_interconnect_0:hdd_avalon_master_address
	wire         hdd_avalon_master_write;                                   // hdd:sd_master_write -> mm_interconnect_0:hdd_avalon_master_write
	wire         hdd_avalon_master_read;                                    // hdd:sd_master_read -> mm_interconnect_0:hdd_avalon_master_read
	wire  [31:0] hdd_avalon_master_readdata;                                // mm_interconnect_0:hdd_avalon_master_readdata -> hdd:sd_master_readdata
	wire         hdd_avalon_master_readdatavalid;                           // mm_interconnect_0:hdd_avalon_master_readdatavalid -> hdd:sd_master_readdatavalid
	wire   [2:0] pc_bus_avalon_sdram_master_burstcount;                     // pc_bus:sdram_burstcount -> mm_interconnect_0:pc_bus_avalon_sdram_master_burstcount
	wire         pc_bus_avalon_sdram_master_waitrequest;                    // mm_interconnect_0:pc_bus_avalon_sdram_master_waitrequest -> pc_bus:sdram_waitrequest
	wire  [31:0] pc_bus_avalon_sdram_master_writedata;                      // pc_bus:sdram_writedata -> mm_interconnect_0:pc_bus_avalon_sdram_master_writedata
	wire  [31:0] pc_bus_avalon_sdram_master_address;                        // pc_bus:sdram_address -> mm_interconnect_0:pc_bus_avalon_sdram_master_address
	wire         pc_bus_avalon_sdram_master_write;                          // pc_bus:sdram_write -> mm_interconnect_0:pc_bus_avalon_sdram_master_write
	wire         pc_bus_avalon_sdram_master_read;                           // pc_bus:sdram_read -> mm_interconnect_0:pc_bus_avalon_sdram_master_read
	wire  [31:0] pc_bus_avalon_sdram_master_readdata;                       // mm_interconnect_0:pc_bus_avalon_sdram_master_readdata -> pc_bus:sdram_readdata
	wire         pc_bus_avalon_sdram_master_readdatavalid;                  // mm_interconnect_0:pc_bus_avalon_sdram_master_readdatavalid -> pc_bus:sdram_readdatavalid
	wire   [3:0] pc_bus_avalon_sdram_master_byteenable;                     // pc_bus:sdram_byteenable -> mm_interconnect_0:pc_bus_avalon_sdram_master_byteenable
	wire         pc_dma_avalon_master_waitrequest;                          // mm_interconnect_0:pc_dma_avalon_master_waitrequest -> pc_dma:avm_waitrequest
	wire   [7:0] pc_dma_avalon_master_writedata;                            // pc_dma:avm_writedata -> mm_interconnect_0:pc_dma_avalon_master_writedata
	wire  [31:0] pc_dma_avalon_master_address;                              // pc_dma:avm_address -> mm_interconnect_0:pc_dma_avalon_master_address
	wire         pc_dma_avalon_master_write;                                // pc_dma:avm_write -> mm_interconnect_0:pc_dma_avalon_master_write
	wire         pc_dma_avalon_master_read;                                 // pc_dma:avm_read -> mm_interconnect_0:pc_dma_avalon_master_read
	wire   [7:0] pc_dma_avalon_master_readdata;                             // mm_interconnect_0:pc_dma_avalon_master_readdata -> pc_dma:avm_readdata
	wire         pc_dma_avalon_master_readdatavalid;                        // mm_interconnect_0:pc_dma_avalon_master_readdatavalid -> pc_dma:avm_readdatavalid
	wire         driver_sd_avalon_master_0_waitrequest;                     // mm_interconnect_0:driver_sd_avalon_master_0_waitrequest -> driver_sd:avm_waitrequest
	wire  [31:0] driver_sd_avalon_master_0_address;                         // driver_sd:avm_address -> mm_interconnect_0:driver_sd_avalon_master_0_address
	wire  [31:0] driver_sd_avalon_master_0_writedata;                       // driver_sd:avm_writedata -> mm_interconnect_0:driver_sd_avalon_master_0_writedata
	wire         driver_sd_avalon_master_0_write;                           // driver_sd:avm_write -> mm_interconnect_0:driver_sd_avalon_master_0_write
	wire         driver_sd_avalon_master_0_read;                            // driver_sd:avm_read -> mm_interconnect_0:driver_sd_avalon_master_0_read
	wire  [31:0] driver_sd_avalon_master_0_readdata;                        // mm_interconnect_0:driver_sd_avalon_master_0_readdata -> driver_sd:avm_readdata
	wire         driver_sd_avalon_master_0_readdatavalid;                   // mm_interconnect_0:driver_sd_avalon_master_0_readdatavalid -> driver_sd:avm_readdatavalid
	wire         nios2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_instruction_master_waitrequest -> nios2:i_waitrequest
	wire  [16:0] nios2_instruction_master_address;                          // nios2:i_address -> mm_interconnect_0:nios2_instruction_master_address
	wire         nios2_instruction_master_read;                             // nios2:i_read -> mm_interconnect_0:nios2_instruction_master_read
	wire  [31:0] nios2_instruction_master_readdata;                         // mm_interconnect_0:nios2_instruction_master_readdata -> nios2:i_readdata
	wire         ao486_avalon_io_waitrequest;                               // mm_interconnect_0:ao486_avalon_io_waitrequest -> ao486:avalon_io_waitrequest
	wire  [31:0] ao486_avalon_io_writedata;                                 // ao486:avalon_io_writedata -> mm_interconnect_0:ao486_avalon_io_writedata
	wire  [15:0] ao486_avalon_io_address;                                   // ao486:avalon_io_address -> mm_interconnect_0:ao486_avalon_io_address
	wire         ao486_avalon_io_write;                                     // ao486:avalon_io_write -> mm_interconnect_0:ao486_avalon_io_write
	wire         ao486_avalon_io_read;                                      // ao486:avalon_io_read -> mm_interconnect_0:ao486_avalon_io_read
	wire  [31:0] ao486_avalon_io_readdata;                                  // mm_interconnect_0:ao486_avalon_io_readdata -> ao486:avalon_io_readdata
	wire         ao486_avalon_io_readdatavalid;                             // mm_interconnect_0:ao486_avalon_io_readdatavalid -> ao486:avalon_io_readdatavalid
	wire   [3:0] ao486_avalon_io_byteenable;                                // ao486:avalon_io_byteenable -> mm_interconnect_0:ao486_avalon_io_byteenable
	wire         mm_interconnect_0_nios2_jtag_debug_module_waitrequest;     // nios2:jtag_debug_module_waitrequest -> mm_interconnect_0:nios2_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_writedata;       // mm_interconnect_0:nios2_jtag_debug_module_writedata -> nios2:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_nios2_jtag_debug_module_address;         // mm_interconnect_0:nios2_jtag_debug_module_address -> nios2:jtag_debug_module_address
	wire         mm_interconnect_0_nios2_jtag_debug_module_write;           // mm_interconnect_0:nios2_jtag_debug_module_write -> nios2:jtag_debug_module_write
	wire         mm_interconnect_0_nios2_jtag_debug_module_read;            // mm_interconnect_0:nios2_jtag_debug_module_read -> nios2:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_nios2_jtag_debug_module_readdata;        // nios2:jtag_debug_module_readdata -> mm_interconnect_0:nios2_jtag_debug_module_readdata
	wire         mm_interconnect_0_nios2_jtag_debug_module_debugaccess;     // mm_interconnect_0:nios2_jtag_debug_module_debugaccess -> nios2:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_nios2_jtag_debug_module_byteenable;      // mm_interconnect_0:nios2_jtag_debug_module_byteenable -> nios2:jtag_debug_module_byteenable
	wire  [31:0] mm_interconnect_0_onchip_for_nios2_s1_writedata;           // mm_interconnect_0:onchip_for_nios2_s1_writedata -> onchip_for_nios2:writedata
	wire  [12:0] mm_interconnect_0_onchip_for_nios2_s1_address;             // mm_interconnect_0:onchip_for_nios2_s1_address -> onchip_for_nios2:address
	wire         mm_interconnect_0_onchip_for_nios2_s1_chipselect;          // mm_interconnect_0:onchip_for_nios2_s1_chipselect -> onchip_for_nios2:chipselect
	wire         mm_interconnect_0_onchip_for_nios2_s1_clken;               // mm_interconnect_0:onchip_for_nios2_s1_clken -> onchip_for_nios2:clken
	wire         mm_interconnect_0_onchip_for_nios2_s1_write;               // mm_interconnect_0:onchip_for_nios2_s1_write -> onchip_for_nios2:write
	wire  [31:0] mm_interconnect_0_onchip_for_nios2_s1_readdata;            // onchip_for_nios2:readdata -> mm_interconnect_0:onchip_for_nios2_s1_readdata
	wire   [3:0] mm_interconnect_0_onchip_for_nios2_s1_byteenable;          // mm_interconnect_0:onchip_for_nios2_s1_byteenable -> onchip_for_nios2:byteenable
	wire  [31:0] mm_interconnect_0_pc_bus_ctrl_writedata;                   // mm_interconnect_0:pc_bus_ctrl_writedata -> pc_bus:ctrl_writedata
	wire   [1:0] mm_interconnect_0_pc_bus_ctrl_address;                     // mm_interconnect_0:pc_bus_ctrl_address -> pc_bus:ctrl_address
	wire         mm_interconnect_0_pc_bus_ctrl_write;                       // mm_interconnect_0:pc_bus_ctrl_write -> pc_bus:ctrl_write
	wire  [31:0] mm_interconnect_0_vga_sys_writedata;                       // mm_interconnect_0:vga_sys_writedata -> vga:sys_writedata
	wire   [7:0] mm_interconnect_0_vga_sys_address;                         // mm_interconnect_0:vga_sys_address -> vga:sys_address
	wire         mm_interconnect_0_vga_sys_write;                           // mm_interconnect_0:vga_sys_write -> vga:sys_write
	wire         mm_interconnect_0_vga_sys_read;                            // mm_interconnect_0:vga_sys_read -> vga:sys_read
	wire  [31:0] mm_interconnect_0_vga_sys_readdata;                        // vga:sys_readdata -> mm_interconnect_0:vga_sys_readdata
	wire  [31:0] mm_interconnect_0_sound_mgmt_writedata;                    // mm_interconnect_0:sound_mgmt_writedata -> sound:mgmt_writedata
	wire   [8:0] mm_interconnect_0_sound_mgmt_address;                      // mm_interconnect_0:sound_mgmt_address -> sound:mgmt_address
	wire         mm_interconnect_0_sound_mgmt_write;                        // mm_interconnect_0:sound_mgmt_write -> sound:mgmt_write
	wire  [31:0] mm_interconnect_0_rtc_mgmt_writedata;                      // mm_interconnect_0:rtc_mgmt_writedata -> rtc:mgmt_writedata
	wire   [7:0] mm_interconnect_0_rtc_mgmt_address;                        // mm_interconnect_0:rtc_mgmt_address -> rtc:mgmt_address
	wire         mm_interconnect_0_rtc_mgmt_write;                          // mm_interconnect_0:rtc_mgmt_write -> rtc:mgmt_write
	wire  [31:0] mm_interconnect_0_pit_mgmt_writedata;                      // mm_interconnect_0:pit_mgmt_writedata -> pit:mgmt_writedata
	wire   [0:0] mm_interconnect_0_pit_mgmt_address;                        // mm_interconnect_0:pit_mgmt_address -> pit:mgmt_address
	wire         mm_interconnect_0_pit_mgmt_write;                          // mm_interconnect_0:pit_mgmt_write -> pit:mgmt_write
	wire  [31:0] mm_interconnect_0_hdd_mgmt_writedata;                      // mm_interconnect_0:hdd_mgmt_writedata -> hdd:mgmt_writedata
	wire   [2:0] mm_interconnect_0_hdd_mgmt_address;                        // mm_interconnect_0:hdd_mgmt_address -> hdd:mgmt_address
	wire         mm_interconnect_0_hdd_mgmt_write;                          // mm_interconnect_0:hdd_mgmt_write -> hdd:mgmt_write
	wire  [31:0] mm_interconnect_0_floppy_mgmt_writedata;                   // mm_interconnect_0:floppy_mgmt_writedata -> floppy:mgmt_writedata
	wire   [3:0] mm_interconnect_0_floppy_mgmt_address;                     // mm_interconnect_0:floppy_mgmt_address -> floppy:mgmt_address
	wire         mm_interconnect_0_floppy_mgmt_write;                       // mm_interconnect_0:floppy_mgmt_write -> floppy:mgmt_write
	wire  [31:0] mm_interconnect_0_pio_input_s1_writedata;                  // mm_interconnect_0:pio_input_s1_writedata -> pio_input:writedata
	wire   [1:0] mm_interconnect_0_pio_input_s1_address;                    // mm_interconnect_0:pio_input_s1_address -> pio_input:address
	wire         mm_interconnect_0_pio_input_s1_chipselect;                 // mm_interconnect_0:pio_input_s1_chipselect -> pio_input:chipselect
	wire         mm_interconnect_0_pio_input_s1_write;                      // mm_interconnect_0:pio_input_s1_write -> pio_input:write_n
	wire  [31:0] mm_interconnect_0_pio_input_s1_readdata;                   // pio_input:readdata -> mm_interconnect_0:pio_input_s1_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire  [31:0] mm_interconnect_0_pio_output_s1_writedata;                 // mm_interconnect_0:pio_output_s1_writedata -> pio_output:writedata
	wire   [1:0] mm_interconnect_0_pio_output_s1_address;                   // mm_interconnect_0:pio_output_s1_address -> pio_output:address
	wire         mm_interconnect_0_pio_output_s1_chipselect;                // mm_interconnect_0:pio_output_s1_chipselect -> pio_output:chipselect
	wire         mm_interconnect_0_pio_output_s1_write;                     // mm_interconnect_0:pio_output_s1_write -> pio_output:write_n
	wire  [31:0] mm_interconnect_0_pio_output_s1_readdata;                  // pio_output:readdata -> mm_interconnect_0:pio_output_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                    // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                      // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                        // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                     // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                          // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                           // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                       // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                  // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                     // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire  [31:0] mm_interconnect_0_driver_sd_avalon_slave_0_writedata;      // mm_interconnect_0:driver_sd_avalon_slave_0_writedata -> driver_sd:avs_writedata
	wire   [1:0] mm_interconnect_0_driver_sd_avalon_slave_0_address;        // mm_interconnect_0:driver_sd_avalon_slave_0_address -> driver_sd:avs_address
	wire         mm_interconnect_0_driver_sd_avalon_slave_0_write;          // mm_interconnect_0:driver_sd_avalon_slave_0_write -> driver_sd:avs_write
	wire         mm_interconnect_0_driver_sd_avalon_slave_0_read;           // mm_interconnect_0:driver_sd_avalon_slave_0_read -> driver_sd:avs_read
	wire  [31:0] mm_interconnect_0_driver_sd_avalon_slave_0_readdata;       // driver_sd:avs_readdata -> mm_interconnect_0:driver_sd_avalon_slave_0_readdata
	wire   [7:0] mm_interconnect_0_floppy_sd_slave_writedata;               // mm_interconnect_0:floppy_sd_slave_writedata -> floppy:sd_slave_writedata
	wire   [8:0] mm_interconnect_0_floppy_sd_slave_address;                 // mm_interconnect_0:floppy_sd_slave_address -> floppy:sd_slave_address
	wire         mm_interconnect_0_floppy_sd_slave_write;                   // mm_interconnect_0:floppy_sd_slave_write -> floppy:sd_slave_write
	wire         mm_interconnect_0_floppy_sd_slave_read;                    // mm_interconnect_0:floppy_sd_slave_read -> floppy:sd_slave_read
	wire   [7:0] mm_interconnect_0_floppy_sd_slave_readdata;                // floppy:sd_slave_readdata -> mm_interconnect_0:floppy_sd_slave_readdata
	wire  [31:0] mm_interconnect_0_hdd_sd_slave_writedata;                  // mm_interconnect_0:hdd_sd_slave_writedata -> hdd:sd_slave_writedata
	wire   [8:0] mm_interconnect_0_hdd_sd_slave_address;                    // mm_interconnect_0:hdd_sd_slave_address -> hdd:sd_slave_address
	wire         mm_interconnect_0_hdd_sd_slave_write;                      // mm_interconnect_0:hdd_sd_slave_write -> hdd:sd_slave_write
	wire         mm_interconnect_0_hdd_sd_slave_read;                       // mm_interconnect_0:hdd_sd_slave_read -> hdd:sd_slave_read
	wire  [31:0] mm_interconnect_0_hdd_sd_slave_readdata;                   // hdd:sd_slave_readdata -> mm_interconnect_0:hdd_sd_slave_readdata
	wire   [7:0] mm_interconnect_0_pc_dma_slave_writedata;                  // mm_interconnect_0:pc_dma_slave_writedata -> pc_dma:slave_writedata
	wire   [3:0] mm_interconnect_0_pc_dma_slave_address;                    // mm_interconnect_0:pc_dma_slave_address -> pc_dma:slave_address
	wire         mm_interconnect_0_pc_dma_slave_write;                      // mm_interconnect_0:pc_dma_slave_write -> pc_dma:slave_write
	wire         mm_interconnect_0_pc_dma_slave_read;                       // mm_interconnect_0:pc_dma_slave_read -> pc_dma:slave_read
	wire   [7:0] mm_interconnect_0_pc_dma_slave_readdata;                   // pc_dma:slave_readdata -> mm_interconnect_0:pc_dma_slave_readdata
	wire   [7:0] mm_interconnect_0_pc_dma_page_writedata;                   // mm_interconnect_0:pc_dma_page_writedata -> pc_dma:page_writedata
	wire   [3:0] mm_interconnect_0_pc_dma_page_address;                     // mm_interconnect_0:pc_dma_page_address -> pc_dma:page_address
	wire         mm_interconnect_0_pc_dma_page_write;                       // mm_interconnect_0:pc_dma_page_write -> pc_dma:page_write
	wire         mm_interconnect_0_pc_dma_page_read;                        // mm_interconnect_0:pc_dma_page_read -> pc_dma:page_read
	wire   [7:0] mm_interconnect_0_pc_dma_page_readdata;                    // pc_dma:page_readdata -> mm_interconnect_0:pc_dma_page_readdata
	wire   [7:0] mm_interconnect_0_pc_dma_master_writedata;                 // mm_interconnect_0:pc_dma_master_writedata -> pc_dma:master_writedata
	wire   [4:0] mm_interconnect_0_pc_dma_master_address;                   // mm_interconnect_0:pc_dma_master_address -> pc_dma:master_address
	wire         mm_interconnect_0_pc_dma_master_write;                     // mm_interconnect_0:pc_dma_master_write -> pc_dma:master_write
	wire         mm_interconnect_0_pc_dma_master_read;                      // mm_interconnect_0:pc_dma_master_read -> pc_dma:master_read
	wire   [7:0] mm_interconnect_0_pc_dma_master_readdata;                  // pc_dma:master_readdata -> mm_interconnect_0:pc_dma_master_readdata
	wire   [7:0] mm_interconnect_0_vga_io_b_writedata;                      // mm_interconnect_0:vga_io_b_writedata -> vga:io_b_writedata
	wire   [3:0] mm_interconnect_0_vga_io_b_address;                        // mm_interconnect_0:vga_io_b_address -> vga:io_b_address
	wire         mm_interconnect_0_vga_io_b_write;                          // mm_interconnect_0:vga_io_b_write -> vga:io_b_write
	wire         mm_interconnect_0_vga_io_b_read;                           // mm_interconnect_0:vga_io_b_read -> vga:io_b_read
	wire   [7:0] mm_interconnect_0_vga_io_b_readdata;                       // vga:io_b_readdata -> mm_interconnect_0:vga_io_b_readdata
	wire   [7:0] mm_interconnect_0_vga_io_c_writedata;                      // mm_interconnect_0:vga_io_c_writedata -> vga:io_c_writedata
	wire   [3:0] mm_interconnect_0_vga_io_c_address;                        // mm_interconnect_0:vga_io_c_address -> vga:io_c_address
	wire         mm_interconnect_0_vga_io_c_write;                          // mm_interconnect_0:vga_io_c_write -> vga:io_c_write
	wire         mm_interconnect_0_vga_io_c_read;                           // mm_interconnect_0:vga_io_c_read -> vga:io_c_read
	wire   [7:0] mm_interconnect_0_vga_io_c_readdata;                       // vga:io_c_readdata -> mm_interconnect_0:vga_io_c_readdata
	wire   [7:0] mm_interconnect_0_vga_io_d_writedata;                      // mm_interconnect_0:vga_io_d_writedata -> vga:io_d_writedata
	wire   [3:0] mm_interconnect_0_vga_io_d_address;                        // mm_interconnect_0:vga_io_d_address -> vga:io_d_address
	wire         mm_interconnect_0_vga_io_d_write;                          // mm_interconnect_0:vga_io_d_write -> vga:io_d_write
	wire         mm_interconnect_0_vga_io_d_read;                           // mm_interconnect_0:vga_io_d_read -> vga:io_d_read
	wire   [7:0] mm_interconnect_0_vga_io_d_readdata;                       // vga:io_d_readdata -> mm_interconnect_0:vga_io_d_readdata
	wire   [7:0] mm_interconnect_0_sound_io_writedata;                      // mm_interconnect_0:sound_io_writedata -> sound:io_writedata
	wire   [3:0] mm_interconnect_0_sound_io_address;                        // mm_interconnect_0:sound_io_address -> sound:io_address
	wire         mm_interconnect_0_sound_io_write;                          // mm_interconnect_0:sound_io_write -> sound:io_write
	wire         mm_interconnect_0_sound_io_read;                           // mm_interconnect_0:sound_io_read -> sound:io_read
	wire   [7:0] mm_interconnect_0_sound_io_readdata;                       // sound:io_readdata -> mm_interconnect_0:sound_io_readdata
	wire   [7:0] mm_interconnect_0_sound_fm_writedata;                      // mm_interconnect_0:sound_fm_writedata -> sound:fm_writedata
	wire   [0:0] mm_interconnect_0_sound_fm_address;                        // mm_interconnect_0:sound_fm_address -> sound:fm_address
	wire         mm_interconnect_0_sound_fm_write;                          // mm_interconnect_0:sound_fm_write -> sound:fm_write
	wire         mm_interconnect_0_sound_fm_read;                           // mm_interconnect_0:sound_fm_read -> sound:fm_read
	wire   [7:0] mm_interconnect_0_sound_fm_readdata;                       // sound:fm_readdata -> mm_interconnect_0:sound_fm_readdata
	wire   [7:0] mm_interconnect_0_rtc_io_writedata;                        // mm_interconnect_0:rtc_io_writedata -> rtc:io_writedata
	wire   [0:0] mm_interconnect_0_rtc_io_address;                          // mm_interconnect_0:rtc_io_address -> rtc:io_address
	wire         mm_interconnect_0_rtc_io_write;                            // mm_interconnect_0:rtc_io_write -> rtc:io_write
	wire         mm_interconnect_0_rtc_io_read;                             // mm_interconnect_0:rtc_io_read -> rtc:io_read
	wire   [7:0] mm_interconnect_0_rtc_io_readdata;                         // rtc:io_readdata -> mm_interconnect_0:rtc_io_readdata
	wire   [7:0] mm_interconnect_0_pit_io_writedata;                        // mm_interconnect_0:pit_io_writedata -> pit:io_writedata
	wire   [1:0] mm_interconnect_0_pit_io_address;                          // mm_interconnect_0:pit_io_address -> pit:io_address
	wire         mm_interconnect_0_pit_io_write;                            // mm_interconnect_0:pit_io_write -> pit:io_write
	wire         mm_interconnect_0_pit_io_read;                             // mm_interconnect_0:pit_io_read -> pit:io_read
	wire   [7:0] mm_interconnect_0_pit_io_readdata;                         // pit:io_readdata -> mm_interconnect_0:pit_io_readdata
	wire   [7:0] mm_interconnect_0_pic_master_writedata;                    // mm_interconnect_0:pic_master_writedata -> pic:master_writedata
	wire   [0:0] mm_interconnect_0_pic_master_address;                      // mm_interconnect_0:pic_master_address -> pic:master_address
	wire         mm_interconnect_0_pic_master_write;                        // mm_interconnect_0:pic_master_write -> pic:master_write
	wire         mm_interconnect_0_pic_master_read;                         // mm_interconnect_0:pic_master_read -> pic:master_read
	wire   [7:0] mm_interconnect_0_pic_master_readdata;                     // pic:master_readdata -> mm_interconnect_0:pic_master_readdata
	wire   [7:0] mm_interconnect_0_pic_slave_writedata;                     // mm_interconnect_0:pic_slave_writedata -> pic:slave_writedata
	wire   [0:0] mm_interconnect_0_pic_slave_address;                       // mm_interconnect_0:pic_slave_address -> pic:slave_address
	wire         mm_interconnect_0_pic_slave_write;                         // mm_interconnect_0:pic_slave_write -> pic:slave_write
	wire         mm_interconnect_0_pic_slave_read;                          // mm_interconnect_0:pic_slave_read -> pic:slave_read
	wire   [7:0] mm_interconnect_0_pic_slave_readdata;                      // pic:slave_readdata -> mm_interconnect_0:pic_slave_readdata
	wire  [31:0] mm_interconnect_0_hdd_io_writedata;                        // mm_interconnect_0:hdd_io_writedata -> hdd:io_writedata
	wire   [0:0] mm_interconnect_0_hdd_io_address;                          // mm_interconnect_0:hdd_io_address -> hdd:io_address
	wire         mm_interconnect_0_hdd_io_write;                            // mm_interconnect_0:hdd_io_write -> hdd:io_write
	wire         mm_interconnect_0_hdd_io_read;                             // mm_interconnect_0:hdd_io_read -> hdd:io_read
	wire  [31:0] mm_interconnect_0_hdd_io_readdata;                         // hdd:io_readdata -> mm_interconnect_0:hdd_io_readdata
	wire   [3:0] mm_interconnect_0_hdd_io_byteenable;                       // mm_interconnect_0:hdd_io_byteenable -> hdd:io_byteenable
	wire   [7:0] mm_interconnect_0_floppy_io_writedata;                     // mm_interconnect_0:floppy_io_writedata -> floppy:io_writedata
	wire   [2:0] mm_interconnect_0_floppy_io_address;                       // mm_interconnect_0:floppy_io_address -> floppy:io_address
	wire         mm_interconnect_0_floppy_io_write;                         // mm_interconnect_0:floppy_io_write -> floppy:io_write
	wire         mm_interconnect_0_floppy_io_read;                          // mm_interconnect_0:floppy_io_read -> floppy:io_read
	wire   [7:0] mm_interconnect_0_floppy_io_readdata;                      // floppy:io_readdata -> mm_interconnect_0:floppy_io_readdata
	wire   [7:0] mm_interconnect_0_ps2_io_writedata;                        // mm_interconnect_0:ps2_io_writedata -> ps2:io_writedata
	wire   [2:0] mm_interconnect_0_ps2_io_address;                          // mm_interconnect_0:ps2_io_address -> ps2:io_address
	wire         mm_interconnect_0_ps2_io_write;                            // mm_interconnect_0:ps2_io_write -> ps2:io_write
	wire         mm_interconnect_0_ps2_io_read;                             // mm_interconnect_0:ps2_io_read -> ps2:io_read
	wire   [7:0] mm_interconnect_0_ps2_io_readdata;                         // ps2:io_readdata -> mm_interconnect_0:ps2_io_readdata
	wire   [7:0] mm_interconnect_0_ps2_sysctl_writedata;                    // mm_interconnect_0:ps2_sysctl_writedata -> ps2:sysctl_writedata
	wire   [3:0] mm_interconnect_0_ps2_sysctl_address;                      // mm_interconnect_0:ps2_sysctl_address -> ps2:sysctl_address
	wire         mm_interconnect_0_ps2_sysctl_write;                        // mm_interconnect_0:ps2_sysctl_write -> ps2:sysctl_write
	wire         mm_interconnect_0_ps2_sysctl_read;                         // mm_interconnect_0:ps2_sysctl_read -> ps2:sysctl_read
	wire   [7:0] mm_interconnect_0_ps2_sysctl_readdata;                     // ps2:sysctl_readdata -> mm_interconnect_0:ps2_sysctl_readdata
	wire   [2:0] pc_bus_avalon_vga_master_burstcount;                       // pc_bus:vga_burstcount -> mm_interconnect_1:pc_bus_avalon_vga_master_burstcount
	wire         pc_bus_avalon_vga_master_waitrequest;                      // mm_interconnect_1:pc_bus_avalon_vga_master_waitrequest -> pc_bus:vga_waitrequest
	wire  [31:0] pc_bus_avalon_vga_master_writedata;                        // pc_bus:vga_writedata -> mm_interconnect_1:pc_bus_avalon_vga_master_writedata
	wire  [31:0] pc_bus_avalon_vga_master_address;                          // pc_bus:vga_address -> mm_interconnect_1:pc_bus_avalon_vga_master_address
	wire         pc_bus_avalon_vga_master_write;                            // pc_bus:vga_write -> mm_interconnect_1:pc_bus_avalon_vga_master_write
	wire         pc_bus_avalon_vga_master_read;                             // pc_bus:vga_read -> mm_interconnect_1:pc_bus_avalon_vga_master_read
	wire  [31:0] pc_bus_avalon_vga_master_readdata;                         // mm_interconnect_1:pc_bus_avalon_vga_master_readdata -> pc_bus:vga_readdata
	wire         pc_bus_avalon_vga_master_readdatavalid;                    // mm_interconnect_1:pc_bus_avalon_vga_master_readdatavalid -> pc_bus:vga_readdatavalid
	wire   [3:0] pc_bus_avalon_vga_master_byteenable;                       // pc_bus:vga_byteenable -> mm_interconnect_1:pc_bus_avalon_vga_master_byteenable
	wire   [7:0] mm_interconnect_1_vga_mem_writedata;                       // mm_interconnect_1:vga_mem_writedata -> vga:mem_writedata
	wire  [16:0] mm_interconnect_1_vga_mem_address;                         // mm_interconnect_1:vga_mem_address -> vga:mem_address
	wire         mm_interconnect_1_vga_mem_write;                           // mm_interconnect_1:vga_mem_write -> vga:mem_write
	wire         mm_interconnect_1_vga_mem_read;                            // mm_interconnect_1:vga_mem_read -> vga:mem_read
	wire   [7:0] mm_interconnect_1_vga_mem_readdata;                        // vga:mem_readdata -> mm_interconnect_1:vga_mem_readdata
	wire         ao486_avalon_memory_waitrequest;                           // mm_interconnect_2:ao486_avalon_memory_waitrequest -> ao486:avm_waitrequest
	wire   [2:0] ao486_avalon_memory_burstcount;                            // ao486:avm_burstcount -> mm_interconnect_2:ao486_avalon_memory_burstcount
	wire  [31:0] ao486_avalon_memory_writedata;                             // ao486:avm_writedata -> mm_interconnect_2:ao486_avalon_memory_writedata
	wire  [31:0] ao486_avalon_memory_address;                               // ao486:avm_address -> mm_interconnect_2:ao486_avalon_memory_address
	wire         ao486_avalon_memory_write;                                 // ao486:avm_write -> mm_interconnect_2:ao486_avalon_memory_write
	wire         ao486_avalon_memory_read;                                  // ao486:avm_read -> mm_interconnect_2:ao486_avalon_memory_read
	wire  [31:0] ao486_avalon_memory_readdata;                              // mm_interconnect_2:ao486_avalon_memory_readdata -> ao486:avm_readdata
	wire         ao486_avalon_memory_readdatavalid;                         // mm_interconnect_2:ao486_avalon_memory_readdatavalid -> ao486:avm_readdatavalid
	wire   [3:0] ao486_avalon_memory_byteenable;                            // ao486:avm_byteenable -> mm_interconnect_2:ao486_avalon_memory_byteenable
	wire         mm_interconnect_2_pc_bus_mem_waitrequest;                  // pc_bus:mem_waitrequest -> mm_interconnect_2:pc_bus_mem_waitrequest
	wire   [2:0] mm_interconnect_2_pc_bus_mem_burstcount;                   // mm_interconnect_2:pc_bus_mem_burstcount -> pc_bus:mem_burstcount
	wire  [31:0] mm_interconnect_2_pc_bus_mem_writedata;                    // mm_interconnect_2:pc_bus_mem_writedata -> pc_bus:mem_writedata
	wire  [29:0] mm_interconnect_2_pc_bus_mem_address;                      // mm_interconnect_2:pc_bus_mem_address -> pc_bus:mem_address
	wire         mm_interconnect_2_pc_bus_mem_write;                        // mm_interconnect_2:pc_bus_mem_write -> pc_bus:mem_write
	wire         mm_interconnect_2_pc_bus_mem_read;                         // mm_interconnect_2:pc_bus_mem_read -> pc_bus:mem_read
	wire  [31:0] mm_interconnect_2_pc_bus_mem_readdata;                     // pc_bus:mem_readdata -> mm_interconnect_2:pc_bus_mem_readdata
	wire         mm_interconnect_2_pc_bus_mem_readdatavalid;                // pc_bus:mem_readdatavalid -> mm_interconnect_2:pc_bus_mem_readdatavalid
	wire   [3:0] mm_interconnect_2_pc_bus_mem_byteenable;                   // mm_interconnect_2:pc_bus_mem_byteenable -> pc_bus:mem_byteenable
	wire         sound_sound_master_waitrequest;                            // mm_interconnect_3:sound_sound_master_waitrequest -> sound:avm_waitrequest
	wire   [2:0] sound_sound_master_address;                                // sound:avm_address -> mm_interconnect_3:sound_sound_master_address
	wire  [31:0] sound_sound_master_writedata;                              // sound:avm_writedata -> mm_interconnect_3:sound_sound_master_writedata
	wire         sound_sound_master_write;                                  // sound:avm_write -> mm_interconnect_3:sound_sound_master_write
	wire  [31:0] mm_interconnect_3_driver_sound_sound_slave_writedata;      // mm_interconnect_3:driver_sound_sound_slave_writedata -> driver_sound:avs_writedata
	wire         mm_interconnect_3_driver_sound_sound_slave_write;          // mm_interconnect_3:driver_sound_sound_slave_write -> driver_sound:avs_write
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_d_irq_irq;                                           // irq_mapper:sender_irq -> nios2:d_irq
	wire         irq_mapper_001_receiver0_irq;                              // pit:irq -> irq_mapper_001:receiver0_irq
	wire         irq_mapper_001_receiver1_irq;                              // rtc:irq -> irq_mapper_001:receiver1_irq
	wire         irq_mapper_001_receiver2_irq;                              // sound:irq -> irq_mapper_001:receiver2_irq
	wire         irq_mapper_001_receiver3_irq;                              // hdd:irq -> irq_mapper_001:receiver3_irq
	wire         irq_mapper_001_receiver4_irq;                              // ps2:irq_mouse -> irq_mapper_001:receiver4_irq
	wire         irq_mapper_001_receiver5_irq;                              // ps2:irq_keyb -> irq_mapper_001:receiver5_irq
	wire         irq_mapper_001_receiver6_irq;                              // floppy:irq -> irq_mapper_001:receiver6_irq
	wire  [15:0] pic_interrupt_receiver_irq;                                // irq_mapper_001:sender_irq -> pic:interrupt_input
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [driver_sd:rst_n, floppy:rst_n, hdd:rst_n, irq_mapper:reset, irq_mapper_001:reset, jtag_uart:rst_n, mm_interconnect_0:nios2_reset_n_reset_bridge_in_reset_reset, mm_interconnect_1:pc_bus_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_2:pc_bus_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_3:sound_reset_sink_reset_bridge_in_reset_reset, nios2:reset_n, onchip_for_nios2:reset, pc_bus:rst_n, pc_dma:rst_n, pic:rst_n, pio_input:reset_n, pio_output:reset_n, pit:rst_n, ps2:rst_n, rst_translator:in_reset, rtc:rst_n, sdram:reset_n, sound:rst_n]
	wire         rst_controller_reset_out_reset_req;                        // rst_controller:reset_req -> [nios2:reset_req, onchip_for_nios2:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [mm_interconnect_0:vga_reset_sink_reset_bridge_in_reset_reset, mm_interconnect_1:vga_reset_sink_reset_bridge_in_reset_reset, vga:rst_n]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [driver_sound:rst_n, mm_interconnect_3:driver_sound_reset_sound_reset_bridge_in_reset_reset]

	ao486 ao486 (
		.clk                     (clk_sys_clk),                            //         clock.clk
		.rst_n                   (~reset_only_ao486_reset_out_reset),      //    reset_sink.reset_n
		.avm_address             (ao486_avalon_memory_address),            // avalon_memory.address
		.avm_writedata           (ao486_avalon_memory_writedata),          //              .writedata
		.avm_byteenable          (ao486_avalon_memory_byteenable),         //              .byteenable
		.avm_burstcount          (ao486_avalon_memory_burstcount),         //              .burstcount
		.avm_write               (ao486_avalon_memory_write),              //              .write
		.avm_read                (ao486_avalon_memory_read),               //              .read
		.avm_waitrequest         (ao486_avalon_memory_waitrequest),        //              .waitrequest
		.avm_readdatavalid       (ao486_avalon_memory_readdatavalid),      //              .readdatavalid
		.avm_readdata            (ao486_avalon_memory_readdata),           //              .readdata
		.interrupt_do            (pic_conduit_interrupt_interrupt_do),     //     interrupt.interrupt_do
		.interrupt_vector        (pic_conduit_interrupt_interrupt_vector), //              .interrupt_vector
		.interrupt_done          (ao486_interrupt_interrupt_done),         //              .interrupt_done
		.avalon_io_address       (ao486_avalon_io_address),                //     avalon_io.address
		.avalon_io_byteenable    (ao486_avalon_io_byteenable),             //              .byteenable
		.avalon_io_read          (ao486_avalon_io_read),                   //              .read
		.avalon_io_readdatavalid (ao486_avalon_io_readdatavalid),          //              .readdatavalid
		.avalon_io_readdata      (ao486_avalon_io_readdata),               //              .readdata
		.avalon_io_write         (ao486_avalon_io_write),                  //              .write
		.avalon_io_writedata     (ao486_avalon_io_writedata),              //              .writedata
		.avalon_io_waitrequest   (ao486_avalon_io_waitrequest)             //              .waitrequest
	);

	system_nios2 nios2 (
		.clk                                   (clk_sys_clk),                                           //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                       //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                    //                          .reset_req
		.d_address                             (nios2_data_master_address),                             //               data_master.address
		.d_byteenable                          (nios2_data_master_byteenable),                          //                          .byteenable
		.d_read                                (nios2_data_master_read),                                //                          .read
		.d_readdata                            (nios2_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (nios2_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (nios2_data_master_write),                               //                          .write
		.d_writedata                           (nios2_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (nios2_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (nios2_instruction_master_address),                      //        instruction_master.address
		.i_read                                (nios2_instruction_master_read),                         //                          .read
		.i_readdata                            (nios2_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (nios2_instruction_master_waitrequest),                  //                          .waitrequest
		.d_irq                                 (nios2_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (nios2_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_nios2_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_nios2_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_nios2_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_nios2_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_nios2_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_nios2_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_nios2_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_nios2_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                       // custom_instruction_master.readra
	);

	system_onchip_for_nios2 onchip_for_nios2 (
		.clk        (clk_sys_clk),                                      //   clk1.clk
		.address    (mm_interconnect_0_onchip_for_nios2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_for_nios2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_for_nios2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_for_nios2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_for_nios2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_for_nios2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_for_nios2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req)                //       .reset_req
	);

	system_jtag_uart jtag_uart (
		.clk            (clk_sys_clk),                                               //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                           //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	pc_bus pc_bus (
		.clk                 (clk_sys_clk),                                //               clock.clk
		.ctrl_address        (mm_interconnect_0_pc_bus_ctrl_address),      //                ctrl.address
		.ctrl_write          (mm_interconnect_0_pc_bus_ctrl_write),        //                    .write
		.ctrl_writedata      (mm_interconnect_0_pc_bus_ctrl_writedata),    //                    .writedata
		.mem_address         (mm_interconnect_2_pc_bus_mem_address),       //                 mem.address
		.mem_byteenable      (mm_interconnect_2_pc_bus_mem_byteenable),    //                    .byteenable
		.mem_read            (mm_interconnect_2_pc_bus_mem_read),          //                    .read
		.mem_readdata        (mm_interconnect_2_pc_bus_mem_readdata),      //                    .readdata
		.mem_write           (mm_interconnect_2_pc_bus_mem_write),         //                    .write
		.mem_writedata       (mm_interconnect_2_pc_bus_mem_writedata),     //                    .writedata
		.mem_waitrequest     (mm_interconnect_2_pc_bus_mem_waitrequest),   //                    .waitrequest
		.mem_readdatavalid   (mm_interconnect_2_pc_bus_mem_readdatavalid), //                    .readdatavalid
		.mem_burstcount      (mm_interconnect_2_pc_bus_mem_burstcount),    //                    .burstcount
		.rst_n               (~rst_controller_reset_out_reset),            //          reset_sink.reset_n
		.vga_address         (pc_bus_avalon_vga_master_address),           //   avalon_vga_master.address
		.vga_byteenable      (pc_bus_avalon_vga_master_byteenable),        //                    .byteenable
		.vga_read            (pc_bus_avalon_vga_master_read),              //                    .read
		.vga_readdata        (pc_bus_avalon_vga_master_readdata),          //                    .readdata
		.vga_write           (pc_bus_avalon_vga_master_write),             //                    .write
		.vga_writedata       (pc_bus_avalon_vga_master_writedata),         //                    .writedata
		.vga_waitrequest     (pc_bus_avalon_vga_master_waitrequest),       //                    .waitrequest
		.vga_readdatavalid   (pc_bus_avalon_vga_master_readdatavalid),     //                    .readdatavalid
		.vga_burstcount      (pc_bus_avalon_vga_master_burstcount),        //                    .burstcount
		.sdram_address       (pc_bus_avalon_sdram_master_address),         // avalon_sdram_master.address
		.sdram_byteenable    (pc_bus_avalon_sdram_master_byteenable),      //                    .byteenable
		.sdram_read          (pc_bus_avalon_sdram_master_read),            //                    .read
		.sdram_readdata      (pc_bus_avalon_sdram_master_readdata),        //                    .readdata
		.sdram_write         (pc_bus_avalon_sdram_master_write),           //                    .write
		.sdram_writedata     (pc_bus_avalon_sdram_master_writedata),       //                    .writedata
		.sdram_waitrequest   (pc_bus_avalon_sdram_master_waitrequest),     //                    .waitrequest
		.sdram_readdatavalid (pc_bus_avalon_sdram_master_readdatavalid),   //                    .readdatavalid
		.sdram_burstcount    (pc_bus_avalon_sdram_master_burstcount)       //                    .burstcount
	);

	vga vga (
		.sys_address    (mm_interconnect_0_vga_sys_address),    //        sys.address
		.sys_read       (mm_interconnect_0_vga_sys_read),       //           .read
		.sys_readdata   (mm_interconnect_0_vga_sys_readdata),   //           .readdata
		.sys_write      (mm_interconnect_0_vga_sys_write),      //           .write
		.sys_writedata  (mm_interconnect_0_vga_sys_writedata),  //           .writedata
		.io_b_address   (mm_interconnect_0_vga_io_b_address),   //       io_b.address
		.io_b_read      (mm_interconnect_0_vga_io_b_read),      //           .read
		.io_b_readdata  (mm_interconnect_0_vga_io_b_readdata),  //           .readdata
		.io_b_write     (mm_interconnect_0_vga_io_b_write),     //           .write
		.io_b_writedata (mm_interconnect_0_vga_io_b_writedata), //           .writedata
		.io_c_address   (mm_interconnect_0_vga_io_c_address),   //       io_c.address
		.io_c_read      (mm_interconnect_0_vga_io_c_read),      //           .read
		.io_c_readdata  (mm_interconnect_0_vga_io_c_readdata),  //           .readdata
		.io_c_write     (mm_interconnect_0_vga_io_c_write),     //           .write
		.io_c_writedata (mm_interconnect_0_vga_io_c_writedata), //           .writedata
		.io_d_address   (mm_interconnect_0_vga_io_d_address),   //       io_d.address
		.io_d_read      (mm_interconnect_0_vga_io_d_read),      //           .read
		.io_d_readdata  (mm_interconnect_0_vga_io_d_readdata),  //           .readdata
		.io_d_write     (mm_interconnect_0_vga_io_d_write),     //           .write
		.io_d_writedata (mm_interconnect_0_vga_io_d_writedata), //           .writedata
		.mem_address    (mm_interconnect_1_vga_mem_address),    //        mem.address
		.mem_read       (mm_interconnect_1_vga_mem_read),       //           .read
		.mem_readdata   (mm_interconnect_1_vga_mem_readdata),   //           .readdata
		.mem_write      (mm_interconnect_1_vga_mem_write),      //           .write
		.mem_writedata  (mm_interconnect_1_vga_mem_writedata),  //           .writedata
		.clk_26         (clk_vga_clk),                          // clock_sink.clk
		.rst_n          (~rst_controller_001_reset_out_reset),  // reset_sink.reset_n
		.vga_clock      (export_vga_clock),                     // export_vga.export
		.vga_sync_n     (export_vga_sync_n),                    //           .export
		.vga_blank_n    (export_vga_blank_n),                   //           .export
		.vga_horiz_sync (export_vga_horiz_sync),                //           .export
		.vga_vert_sync  (export_vga_vert_sync),                 //           .export
		.vga_r          (export_vga_r),                         //           .export
		.vga_g          (export_vga_g),                         //           .export
		.vga_b          (export_vga_b)                          //           .export
	);

	system_sdram sdram (
		.clk            (clk_sys_clk),                              //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_conduit_end_addr),                   //  wire.export
		.zs_ba          (sdram_conduit_end_ba),                     //      .export
		.zs_cas_n       (sdram_conduit_end_cas_n),                  //      .export
		.zs_cke         (sdram_conduit_end_cke),                    //      .export
		.zs_cs_n        (sdram_conduit_end_cs_n),                   //      .export
		.zs_dq          (sdram_conduit_end_dq),                     //      .export
		.zs_dqm         (sdram_conduit_end_dqm),                    //      .export
		.zs_ras_n       (sdram_conduit_end_ras_n),                  //      .export
		.zs_we_n        (sdram_conduit_end_we_n)                    //      .export
	);

	sound sound (
		.clk                        (clk_sys_clk),                              //                    clock.clk
		.io_address                 (mm_interconnect_0_sound_io_address),       //                       io.address
		.io_read                    (mm_interconnect_0_sound_io_read),          //                         .read
		.io_readdata                (mm_interconnect_0_sound_io_readdata),      //                         .readdata
		.io_write                   (mm_interconnect_0_sound_io_write),         //                         .write
		.io_writedata               (mm_interconnect_0_sound_io_writedata),     //                         .writedata
		.fm_address                 (mm_interconnect_0_sound_fm_address),       //                       fm.address
		.fm_read                    (mm_interconnect_0_sound_fm_read),          //                         .read
		.fm_readdata                (mm_interconnect_0_sound_fm_readdata),      //                         .readdata
		.fm_write                   (mm_interconnect_0_sound_fm_write),         //                         .write
		.fm_writedata               (mm_interconnect_0_sound_fm_writedata),     //                         .writedata
		.mgmt_address               (mm_interconnect_0_sound_mgmt_address),     //                     mgmt.address
		.mgmt_write                 (mm_interconnect_0_sound_mgmt_write),       //                         .write
		.mgmt_writedata             (mm_interconnect_0_sound_mgmt_writedata),   //                         .writedata
		.rst_n                      (~rst_controller_reset_out_reset),          //               reset_sink.reset_n
		.irq                        (irq_mapper_001_receiver2_irq),             //         interrupt_sender.irq
		.avm_write                  (sound_sound_master_write),                 //             sound_master.write
		.avm_writedata              (sound_sound_master_writedata),             //                         .writedata
		.avm_address                (sound_sound_master_address),               //                         .address
		.avm_waitrequest            (sound_sound_master_waitrequest),           //                         .waitrequest
		.speaker_enable             (pit_conduit_speaker_enable),               //          conduit_speaker.export
		.speaker_out                (pit_conduit_speaker_out),                  //                         .export
		.dma_soundblaster_req       (sound_conduit_dma_soundblaster_req),       // conduit_dma_soundblaster.export
		.dma_soundblaster_ack       (pc_dma_conduit_dma_soundblaster_ack),      //                         .export
		.dma_soundblaster_terminal  (pc_dma_conduit_dma_soundblaster_terminal), //                         .export
		.dma_soundblaster_readdata  (pc_dma_conduit_dma_soundblaster_readdata), //                         .export
		.dma_soundblaster_writedata (sound_conduit_dma_soundblaster_writedata)  //                         .export
	);

	rtc rtc (
		.clk            (clk_sys_clk),                          //         clock.clk
		.io_address     (mm_interconnect_0_rtc_io_address),     //            io.address
		.io_read        (mm_interconnect_0_rtc_io_read),        //              .read
		.io_readdata    (mm_interconnect_0_rtc_io_readdata),    //              .readdata
		.io_write       (mm_interconnect_0_rtc_io_write),       //              .write
		.io_writedata   (mm_interconnect_0_rtc_io_writedata),   //              .writedata
		.mgmt_address   (mm_interconnect_0_rtc_mgmt_address),   //          mgmt.address
		.mgmt_write     (mm_interconnect_0_rtc_mgmt_write),     //              .write
		.mgmt_writedata (mm_interconnect_0_rtc_mgmt_writedata), //              .writedata
		.rst_n          (~rst_controller_reset_out_reset),      //    reset_sink.reset_n
		.irq            (irq_mapper_001_receiver1_irq)          // interrupt_rtc.irq
	);

	pit pit (
		.clk                   (clk_sys_clk),                          //               clock.clk
		.io_address            (mm_interconnect_0_pit_io_address),     //                  io.address
		.io_read               (mm_interconnect_0_pit_io_read),        //                    .read
		.io_readdata           (mm_interconnect_0_pit_io_readdata),    //                    .readdata
		.io_write              (mm_interconnect_0_pit_io_write),       //                    .write
		.io_writedata          (mm_interconnect_0_pit_io_writedata),   //                    .writedata
		.mgmt_address          (mm_interconnect_0_pit_mgmt_address),   //                mgmt.address
		.mgmt_write            (mm_interconnect_0_pit_mgmt_write),     //                    .write
		.mgmt_writedata        (mm_interconnect_0_pit_mgmt_writedata), //                    .writedata
		.rst_n                 (~rst_controller_reset_out_reset),      //          reset_sink.reset_n
		.speaker_61h_read      (ps2_conduit_speaker_61h_read),         // conduit_speaker_61h.export
		.speaker_61h_readdata  (pit_conduit_speaker_61h_readdata),     //                    .export
		.speaker_61h_write     (ps2_conduit_speaker_61h_write),        //                    .export
		.speaker_61h_writedata (ps2_conduit_speaker_61h_writedata),    //                    .export
		.speaker_enable        (pit_conduit_speaker_enable),           //     conduit_speaker.export
		.speaker_out           (pit_conduit_speaker_out),              //                    .export
		.irq                   (irq_mapper_001_receiver0_irq)          //       interrupt_pit.irq
	);

	pic pic (
		.clk              (clk_sys_clk),                            //              clock.clk
		.master_address   (mm_interconnect_0_pic_master_address),   //             master.address
		.master_read      (mm_interconnect_0_pic_master_read),      //                   .read
		.master_readdata  (mm_interconnect_0_pic_master_readdata),  //                   .readdata
		.master_write     (mm_interconnect_0_pic_master_write),     //                   .write
		.master_writedata (mm_interconnect_0_pic_master_writedata), //                   .writedata
		.slave_address    (mm_interconnect_0_pic_slave_address),    //              slave.address
		.slave_read       (mm_interconnect_0_pic_slave_read),       //                   .read
		.slave_readdata   (mm_interconnect_0_pic_slave_readdata),   //                   .readdata
		.slave_write      (mm_interconnect_0_pic_slave_write),      //                   .write
		.slave_writedata  (mm_interconnect_0_pic_slave_writedata),  //                   .writedata
		.rst_n            (~rst_controller_reset_out_reset),        //         reset_sink.reset_n
		.interrupt_vector (pic_conduit_interrupt_interrupt_vector), //  conduit_interrupt.interrupt_vector
		.interrupt_done   (ao486_interrupt_interrupt_done),         //                   .interrupt_done
		.interrupt_do     (pic_conduit_interrupt_interrupt_do),     //                   .interrupt_do
		.interrupt_input  (pic_interrupt_receiver_irq)              // interrupt_receiver.irq
	);

	hdd hdd (
		.clk                     (clk_sys_clk),                              //            clock.clk
		.io_address              (mm_interconnect_0_hdd_io_address),         //               io.address
		.io_byteenable           (mm_interconnect_0_hdd_io_byteenable),      //                 .byteenable
		.io_read                 (mm_interconnect_0_hdd_io_read),            //                 .read
		.io_readdata             (mm_interconnect_0_hdd_io_readdata),        //                 .readdata
		.io_write                (mm_interconnect_0_hdd_io_write),           //                 .write
		.io_writedata            (mm_interconnect_0_hdd_io_writedata),       //                 .writedata
		.sd_slave_address        (mm_interconnect_0_hdd_sd_slave_address),   //         sd_slave.address
		.sd_slave_read           (mm_interconnect_0_hdd_sd_slave_read),      //                 .read
		.sd_slave_readdata       (mm_interconnect_0_hdd_sd_slave_readdata),  //                 .readdata
		.sd_slave_write          (mm_interconnect_0_hdd_sd_slave_write),     //                 .write
		.sd_slave_writedata      (mm_interconnect_0_hdd_sd_slave_writedata), //                 .writedata
		.mgmt_address            (mm_interconnect_0_hdd_mgmt_address),       //             mgmt.address
		.mgmt_write              (mm_interconnect_0_hdd_mgmt_write),         //                 .write
		.mgmt_writedata          (mm_interconnect_0_hdd_mgmt_writedata),     //                 .writedata
		.rst_n                   (~rst_controller_reset_out_reset),          //       reset_sink.reset_n
		.irq                     (irq_mapper_001_receiver3_irq),             // interrupt_sender.irq
		.sd_master_address       (hdd_avalon_master_address),                //    avalon_master.address
		.sd_master_waitrequest   (hdd_avalon_master_waitrequest),            //                 .waitrequest
		.sd_master_read          (hdd_avalon_master_read),                   //                 .read
		.sd_master_readdatavalid (hdd_avalon_master_readdatavalid),          //                 .readdatavalid
		.sd_master_readdata      (hdd_avalon_master_readdata),               //                 .readdata
		.sd_master_write         (hdd_avalon_master_write),                  //                 .write
		.sd_master_writedata     (hdd_avalon_master_writedata),              //                 .writedata
		.ide_3f6_read            (floppy_conduit_ide_3f6_read),              //  conduit_ide_3f6.export
		.ide_3f6_readdata        (hdd_conduit_ide_3f6_readdata),             //                 .export
		.ide_3f6_write           (floppy_conduit_ide_3f6_write),             //                 .export
		.ide_3f6_writedata       (floppy_conduit_ide_3f6_writedata)          //                 .export
	);

	floppy floppy (
		.clk                     (clk_sys_clk),                                 //              clock.clk
		.io_address              (mm_interconnect_0_floppy_io_address),         //                 io.address
		.io_read                 (mm_interconnect_0_floppy_io_read),            //                   .read
		.io_readdata             (mm_interconnect_0_floppy_io_readdata),        //                   .readdata
		.io_write                (mm_interconnect_0_floppy_io_write),           //                   .write
		.io_writedata            (mm_interconnect_0_floppy_io_writedata),       //                   .writedata
		.sd_slave_address        (mm_interconnect_0_floppy_sd_slave_address),   //           sd_slave.address
		.sd_slave_read           (mm_interconnect_0_floppy_sd_slave_read),      //                   .read
		.sd_slave_readdata       (mm_interconnect_0_floppy_sd_slave_readdata),  //                   .readdata
		.sd_slave_write          (mm_interconnect_0_floppy_sd_slave_write),     //                   .write
		.sd_slave_writedata      (mm_interconnect_0_floppy_sd_slave_writedata), //                   .writedata
		.mgmt_address            (mm_interconnect_0_floppy_mgmt_address),       //               mgmt.address
		.mgmt_write              (mm_interconnect_0_floppy_mgmt_write),         //                   .write
		.mgmt_writedata          (mm_interconnect_0_floppy_mgmt_writedata),     //                   .writedata
		.rst_n                   (~rst_controller_reset_out_reset),             //         reset_sink.reset_n
		.sd_master_address       (floppy_avalon_master_address),                //      avalon_master.address
		.sd_master_waitrequest   (floppy_avalon_master_waitrequest),            //                   .waitrequest
		.sd_master_read          (floppy_avalon_master_read),                   //                   .read
		.sd_master_readdatavalid (floppy_avalon_master_readdatavalid),          //                   .readdatavalid
		.sd_master_readdata      (floppy_avalon_master_readdata),               //                   .readdata
		.sd_master_write         (floppy_avalon_master_write),                  //                   .write
		.sd_master_writedata     (floppy_avalon_master_writedata),              //                   .writedata
		.dma_floppy_req          (floppy_conduit_dma_floppy_req),               // conduit_dma_floppy.export
		.dma_floppy_ack          (pc_dma_conduit_dma_floppy_ack),               //                   .export
		.dma_floppy_terminal     (pc_dma_conduit_dma_floppy_terminal),          //                   .export
		.dma_floppy_readdata     (pc_dma_conduit_dma_floppy_readdata),          //                   .export
		.dma_floppy_writedata    (floppy_conduit_dma_floppy_writedata),         //                   .export
		.ide_3f6_read            (floppy_conduit_ide_3f6_read),                 //    conduit_ide_3f6.export
		.ide_3f6_readdata        (hdd_conduit_ide_3f6_readdata),                //                   .export
		.ide_3f6_write           (floppy_conduit_ide_3f6_write),                //                   .export
		.ide_3f6_writedata       (floppy_conduit_ide_3f6_writedata),            //                   .export
		.irq                     (irq_mapper_001_receiver6_irq)                 //   interrupt_sender.irq
	);

	pc_dma pc_dma (
		.clk                        (clk_sys_clk),                               //                    clock.clk
		.slave_address              (mm_interconnect_0_pc_dma_slave_address),    //                    slave.address
		.slave_read                 (mm_interconnect_0_pc_dma_slave_read),       //                         .read
		.slave_readdata             (mm_interconnect_0_pc_dma_slave_readdata),   //                         .readdata
		.slave_write                (mm_interconnect_0_pc_dma_slave_write),      //                         .write
		.slave_writedata            (mm_interconnect_0_pc_dma_slave_writedata),  //                         .writedata
		.page_address               (mm_interconnect_0_pc_dma_page_address),     //                     page.address
		.page_read                  (mm_interconnect_0_pc_dma_page_read),        //                         .read
		.page_readdata              (mm_interconnect_0_pc_dma_page_readdata),    //                         .readdata
		.page_write                 (mm_interconnect_0_pc_dma_page_write),       //                         .write
		.page_writedata             (mm_interconnect_0_pc_dma_page_writedata),   //                         .writedata
		.master_address             (mm_interconnect_0_pc_dma_master_address),   //                   master.address
		.master_read                (mm_interconnect_0_pc_dma_master_read),      //                         .read
		.master_readdata            (mm_interconnect_0_pc_dma_master_readdata),  //                         .readdata
		.master_write               (mm_interconnect_0_pc_dma_master_write),     //                         .write
		.master_writedata           (mm_interconnect_0_pc_dma_master_writedata), //                         .writedata
		.rst_n                      (~rst_controller_reset_out_reset),           //               reset_sink.reset_n
		.avm_address                (pc_dma_avalon_master_address),              //            avalon_master.address
		.avm_waitrequest            (pc_dma_avalon_master_waitrequest),          //                         .waitrequest
		.avm_read                   (pc_dma_avalon_master_read),                 //                         .read
		.avm_readdatavalid          (pc_dma_avalon_master_readdatavalid),        //                         .readdatavalid
		.avm_readdata               (pc_dma_avalon_master_readdata),             //                         .readdata
		.avm_write                  (pc_dma_avalon_master_write),                //                         .write
		.avm_writedata              (pc_dma_avalon_master_writedata),            //                         .writedata
		.dma_floppy_req             (floppy_conduit_dma_floppy_req),             //       conduit_dma_floppy.export
		.dma_floppy_ack             (pc_dma_conduit_dma_floppy_ack),             //                         .export
		.dma_floppy_terminal        (pc_dma_conduit_dma_floppy_terminal),        //                         .export
		.dma_floppy_readdata        (pc_dma_conduit_dma_floppy_readdata),        //                         .export
		.dma_floppy_writedata       (floppy_conduit_dma_floppy_writedata),       //                         .export
		.dma_soundblaster_req       (sound_conduit_dma_soundblaster_req),        // conduit_dma_soundblaster.export
		.dma_soundblaster_ack       (pc_dma_conduit_dma_soundblaster_ack),       //                         .export
		.dma_soundblaster_terminal  (pc_dma_conduit_dma_soundblaster_terminal),  //                         .export
		.dma_soundblaster_readdata  (pc_dma_conduit_dma_soundblaster_readdata),  //                         .export
		.dma_soundblaster_writedata (sound_conduit_dma_soundblaster_writedata)   //                         .export
	);

	system_pio_input pio_input (
		.clk        (clk_sys_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_pio_input_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_input_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_input_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_input_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_input_s1_readdata),   //                    .readdata
		.in_port    (pio_input_export)                           // external_connection.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_only_ao486 (
		.reset_in0      (reset_only_ao486_reset),           // reset_in0.reset
		.reset_in1      (reset_sys_reset_out_reset),        // reset_in1.reset
		.clk            (clk_sys_clk),                      //       clk.clk
		.reset_out      (reset_only_ao486_reset_out_reset), // reset_out.reset
		.reset_req      (),                                 // (terminated)
		.reset_req_in0  (1'b0),                             // (terminated)
		.reset_req_in1  (1'b0),                             // (terminated)
		.reset_in2      (1'b0),                             // (terminated)
		.reset_req_in2  (1'b0),                             // (terminated)
		.reset_in3      (1'b0),                             // (terminated)
		.reset_req_in3  (1'b0),                             // (terminated)
		.reset_in4      (1'b0),                             // (terminated)
		.reset_req_in4  (1'b0),                             // (terminated)
		.reset_in5      (1'b0),                             // (terminated)
		.reset_req_in5  (1'b0),                             // (terminated)
		.reset_in6      (1'b0),                             // (terminated)
		.reset_req_in6  (1'b0),                             // (terminated)
		.reset_in7      (1'b0),                             // (terminated)
		.reset_req_in7  (1'b0),                             // (terminated)
		.reset_in8      (1'b0),                             // (terminated)
		.reset_req_in8  (1'b0),                             // (terminated)
		.reset_in9      (1'b0),                             // (terminated)
		.reset_req_in9  (1'b0),                             // (terminated)
		.reset_in10     (1'b0),                             // (terminated)
		.reset_req_in10 (1'b0),                             // (terminated)
		.reset_in11     (1'b0),                             // (terminated)
		.reset_req_in11 (1'b0),                             // (terminated)
		.reset_in12     (1'b0),                             // (terminated)
		.reset_req_in12 (1'b0),                             // (terminated)
		.reset_in13     (1'b0),                             // (terminated)
		.reset_req_in13 (1'b0),                             // (terminated)
		.reset_in14     (1'b0),                             // (terminated)
		.reset_req_in14 (1'b0),                             // (terminated)
		.reset_in15     (1'b0),                             // (terminated)
		.reset_req_in15 (1'b0)                              // (terminated)
	);

	system_pio_output pio_output (
		.clk        (clk_sys_clk),                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address    (mm_interconnect_0_pio_output_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_output_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_output_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_output_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_output_s1_readdata),   //                    .readdata
		.out_port   (pio_output_export)                           // external_connection.export
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) reset_sys (
		.reset_in0      (~reset_sys_reset_n),                  // reset_in0.reset
		.reset_in1      (nios2_jtag_debug_module_reset_reset), // reset_in1.reset
		.clk            (clk_sys_clk),                         //       clk.clk
		.reset_out      (reset_sys_reset_out_reset),           // reset_out.reset
		.reset_req      (),                                    // (terminated)
		.reset_req_in0  (1'b0),                                // (terminated)
		.reset_req_in1  (1'b0),                                // (terminated)
		.reset_in2      (1'b0),                                // (terminated)
		.reset_req_in2  (1'b0),                                // (terminated)
		.reset_in3      (1'b0),                                // (terminated)
		.reset_req_in3  (1'b0),                                // (terminated)
		.reset_in4      (1'b0),                                // (terminated)
		.reset_req_in4  (1'b0),                                // (terminated)
		.reset_in5      (1'b0),                                // (terminated)
		.reset_req_in5  (1'b0),                                // (terminated)
		.reset_in6      (1'b0),                                // (terminated)
		.reset_req_in6  (1'b0),                                // (terminated)
		.reset_in7      (1'b0),                                // (terminated)
		.reset_req_in7  (1'b0),                                // (terminated)
		.reset_in8      (1'b0),                                // (terminated)
		.reset_req_in8  (1'b0),                                // (terminated)
		.reset_in9      (1'b0),                                // (terminated)
		.reset_req_in9  (1'b0),                                // (terminated)
		.reset_in10     (1'b0),                                // (terminated)
		.reset_req_in10 (1'b0),                                // (terminated)
		.reset_in11     (1'b0),                                // (terminated)
		.reset_req_in11 (1'b0),                                // (terminated)
		.reset_in12     (1'b0),                                // (terminated)
		.reset_req_in12 (1'b0),                                // (terminated)
		.reset_in13     (1'b0),                                // (terminated)
		.reset_req_in13 (1'b0),                                // (terminated)
		.reset_in14     (1'b0),                                // (terminated)
		.reset_req_in14 (1'b0),                                // (terminated)
		.reset_in15     (1'b0),                                // (terminated)
		.reset_req_in15 (1'b0)                                 // (terminated)
	);

	driver_sound driver_sound (
		.avs_writedata (mm_interconnect_3_driver_sound_sound_slave_writedata), //  sound_slave.writedata
		.avs_write     (mm_interconnect_3_driver_sound_sound_slave_write),     //             .write
		.clk_12        (clk_sound_clk),                                        //  clock_sound.clk
		.rst_n         (~rst_controller_002_reset_out_reset),                  //  reset_sound.reset_n
		.ac_sclk       (export_sound_sclk),                                    // export_sound.export
		.ac_sdat       (export_sound_sdat),                                    //             .export
		.ac_xclk       (export_sound_xclk),                                    //             .export
		.ac_bclk       (export_sound_bclk),                                    //             .export
		.ac_dat        (export_sound_dat),                                     //             .export
		.ac_lr         (export_sound_lr)                                       //             .export
	);

	ps2 ps2 (
		.clk                   (clk_sys_clk),                            //               clock.clk
		.io_address            (mm_interconnect_0_ps2_io_address),       //                  io.address
		.io_read               (mm_interconnect_0_ps2_io_read),          //                    .read
		.io_readdata           (mm_interconnect_0_ps2_io_readdata),      //                    .readdata
		.io_write              (mm_interconnect_0_ps2_io_write),         //                    .write
		.io_writedata          (mm_interconnect_0_ps2_io_writedata),     //                    .writedata
		.sysctl_address        (mm_interconnect_0_ps2_sysctl_address),   //              sysctl.address
		.sysctl_read           (mm_interconnect_0_ps2_sysctl_read),      //                    .read
		.sysctl_readdata       (mm_interconnect_0_ps2_sysctl_readdata),  //                    .readdata
		.sysctl_write          (mm_interconnect_0_ps2_sysctl_write),     //                    .write
		.sysctl_writedata      (mm_interconnect_0_ps2_sysctl_writedata), //                    .writedata
		.rst_n                 (~rst_controller_reset_out_reset),        //          reset_sink.reset_n
		.irq_mouse             (irq_mapper_001_receiver4_irq),           //           irq_mouse.irq
		.ps2_kbclk             (export_ps2_kbclk),                       //          export_ps2.export
		.ps2_kbdat             (export_ps2_kbdat),                       //                    .export
		.ps2_mouseclk          (export_ps2_mouseclk),                    //                    .export
		.ps2_mousedat          (export_ps2_mousedat),                    //                    .export
		.irq_keyb              (irq_mapper_001_receiver5_irq),           //            irq_keyb.irq
		.speaker_61h_read      (ps2_conduit_speaker_61h_read),           // conduit_speaker_61h.export
		.speaker_61h_readdata  (pit_conduit_speaker_61h_readdata),       //                    .export
		.speaker_61h_write     (ps2_conduit_speaker_61h_write),          //                    .export
		.speaker_61h_writedata (ps2_conduit_speaker_61h_writedata),      //                    .export
		.output_a20_enable     (export_ps2_out_port_a20_enable),         // export_ps2_out_port.export
		.output_reset_n        (export_ps2_out_port_reset_n)             //                    .export
	);

	driver_sd driver_sd (
		.clk               (clk_sys_clk),                                          //           clock.clk
		.avs_address       (mm_interconnect_0_driver_sd_avalon_slave_0_address),   //  avalon_slave_0.address
		.avs_read          (mm_interconnect_0_driver_sd_avalon_slave_0_read),      //                .read
		.avs_readdata      (mm_interconnect_0_driver_sd_avalon_slave_0_readdata),  //                .readdata
		.avs_write         (mm_interconnect_0_driver_sd_avalon_slave_0_write),     //                .write
		.avs_writedata     (mm_interconnect_0_driver_sd_avalon_slave_0_writedata), //                .writedata
		.avm_waitrequest   (driver_sd_avalon_master_0_waitrequest),                // avalon_master_0.waitrequest
		.avm_read          (driver_sd_avalon_master_0_read),                       //                .read
		.avm_readdata      (driver_sd_avalon_master_0_readdata),                   //                .readdata
		.avm_readdatavalid (driver_sd_avalon_master_0_readdatavalid),              //                .readdatavalid
		.avm_write         (driver_sd_avalon_master_0_write),                      //                .write
		.avm_writedata     (driver_sd_avalon_master_0_writedata),                  //                .writedata
		.avm_address       (driver_sd_avalon_master_0_address),                    //                .address
		.rst_n             (~rst_controller_reset_out_reset),                      //      reset_sink.reset_n
		.sd_cmd            (sd_cmd_export),                                        //     conduit_cmd.export
		.sd_dat            (sd_dat_export),                                        //     conduit_dat.export
		.sd_clk            (sd_clk_export)                                         //     conduit_clk.export
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clk_sys_clk_clk                              (clk_sys_clk),                                               //                            clk_sys_clk.clk
		.clk_vga_clk_clk                              (clk_vga_clk),                                               //                            clk_vga_clk.clk
		.ao486_reset_sink_reset_bridge_in_reset_reset (reset_only_ao486_reset_out_reset),                          // ao486_reset_sink_reset_bridge_in_reset.reset
		.nios2_reset_n_reset_bridge_in_reset_reset    (rst_controller_reset_out_reset),                            //    nios2_reset_n_reset_bridge_in_reset.reset
		.vga_reset_sink_reset_bridge_in_reset_reset   (rst_controller_001_reset_out_reset),                        //   vga_reset_sink_reset_bridge_in_reset.reset
		.ao486_avalon_io_address                      (ao486_avalon_io_address),                                   //                        ao486_avalon_io.address
		.ao486_avalon_io_waitrequest                  (ao486_avalon_io_waitrequest),                               //                                       .waitrequest
		.ao486_avalon_io_byteenable                   (ao486_avalon_io_byteenable),                                //                                       .byteenable
		.ao486_avalon_io_read                         (ao486_avalon_io_read),                                      //                                       .read
		.ao486_avalon_io_readdata                     (ao486_avalon_io_readdata),                                  //                                       .readdata
		.ao486_avalon_io_readdatavalid                (ao486_avalon_io_readdatavalid),                             //                                       .readdatavalid
		.ao486_avalon_io_write                        (ao486_avalon_io_write),                                     //                                       .write
		.ao486_avalon_io_writedata                    (ao486_avalon_io_writedata),                                 //                                       .writedata
		.driver_sd_avalon_master_0_address            (driver_sd_avalon_master_0_address),                         //              driver_sd_avalon_master_0.address
		.driver_sd_avalon_master_0_waitrequest        (driver_sd_avalon_master_0_waitrequest),                     //                                       .waitrequest
		.driver_sd_avalon_master_0_read               (driver_sd_avalon_master_0_read),                            //                                       .read
		.driver_sd_avalon_master_0_readdata           (driver_sd_avalon_master_0_readdata),                        //                                       .readdata
		.driver_sd_avalon_master_0_readdatavalid      (driver_sd_avalon_master_0_readdatavalid),                   //                                       .readdatavalid
		.driver_sd_avalon_master_0_write              (driver_sd_avalon_master_0_write),                           //                                       .write
		.driver_sd_avalon_master_0_writedata          (driver_sd_avalon_master_0_writedata),                       //                                       .writedata
		.floppy_avalon_master_address                 (floppy_avalon_master_address),                              //                   floppy_avalon_master.address
		.floppy_avalon_master_waitrequest             (floppy_avalon_master_waitrequest),                          //                                       .waitrequest
		.floppy_avalon_master_read                    (floppy_avalon_master_read),                                 //                                       .read
		.floppy_avalon_master_readdata                (floppy_avalon_master_readdata),                             //                                       .readdata
		.floppy_avalon_master_readdatavalid           (floppy_avalon_master_readdatavalid),                        //                                       .readdatavalid
		.floppy_avalon_master_write                   (floppy_avalon_master_write),                                //                                       .write
		.floppy_avalon_master_writedata               (floppy_avalon_master_writedata),                            //                                       .writedata
		.hdd_avalon_master_address                    (hdd_avalon_master_address),                                 //                      hdd_avalon_master.address
		.hdd_avalon_master_waitrequest                (hdd_avalon_master_waitrequest),                             //                                       .waitrequest
		.hdd_avalon_master_read                       (hdd_avalon_master_read),                                    //                                       .read
		.hdd_avalon_master_readdata                   (hdd_avalon_master_readdata),                                //                                       .readdata
		.hdd_avalon_master_readdatavalid              (hdd_avalon_master_readdatavalid),                           //                                       .readdatavalid
		.hdd_avalon_master_write                      (hdd_avalon_master_write),                                   //                                       .write
		.hdd_avalon_master_writedata                  (hdd_avalon_master_writedata),                               //                                       .writedata
		.nios2_data_master_address                    (nios2_data_master_address),                                 //                      nios2_data_master.address
		.nios2_data_master_waitrequest                (nios2_data_master_waitrequest),                             //                                       .waitrequest
		.nios2_data_master_byteenable                 (nios2_data_master_byteenable),                              //                                       .byteenable
		.nios2_data_master_read                       (nios2_data_master_read),                                    //                                       .read
		.nios2_data_master_readdata                   (nios2_data_master_readdata),                                //                                       .readdata
		.nios2_data_master_write                      (nios2_data_master_write),                                   //                                       .write
		.nios2_data_master_writedata                  (nios2_data_master_writedata),                               //                                       .writedata
		.nios2_data_master_debugaccess                (nios2_data_master_debugaccess),                             //                                       .debugaccess
		.nios2_instruction_master_address             (nios2_instruction_master_address),                          //               nios2_instruction_master.address
		.nios2_instruction_master_waitrequest         (nios2_instruction_master_waitrequest),                      //                                       .waitrequest
		.nios2_instruction_master_read                (nios2_instruction_master_read),                             //                                       .read
		.nios2_instruction_master_readdata            (nios2_instruction_master_readdata),                         //                                       .readdata
		.pc_bus_avalon_sdram_master_address           (pc_bus_avalon_sdram_master_address),                        //             pc_bus_avalon_sdram_master.address
		.pc_bus_avalon_sdram_master_waitrequest       (pc_bus_avalon_sdram_master_waitrequest),                    //                                       .waitrequest
		.pc_bus_avalon_sdram_master_burstcount        (pc_bus_avalon_sdram_master_burstcount),                     //                                       .burstcount
		.pc_bus_avalon_sdram_master_byteenable        (pc_bus_avalon_sdram_master_byteenable),                     //                                       .byteenable
		.pc_bus_avalon_sdram_master_read              (pc_bus_avalon_sdram_master_read),                           //                                       .read
		.pc_bus_avalon_sdram_master_readdata          (pc_bus_avalon_sdram_master_readdata),                       //                                       .readdata
		.pc_bus_avalon_sdram_master_readdatavalid     (pc_bus_avalon_sdram_master_readdatavalid),                  //                                       .readdatavalid
		.pc_bus_avalon_sdram_master_write             (pc_bus_avalon_sdram_master_write),                          //                                       .write
		.pc_bus_avalon_sdram_master_writedata         (pc_bus_avalon_sdram_master_writedata),                      //                                       .writedata
		.pc_dma_avalon_master_address                 (pc_dma_avalon_master_address),                              //                   pc_dma_avalon_master.address
		.pc_dma_avalon_master_waitrequest             (pc_dma_avalon_master_waitrequest),                          //                                       .waitrequest
		.pc_dma_avalon_master_read                    (pc_dma_avalon_master_read),                                 //                                       .read
		.pc_dma_avalon_master_readdata                (pc_dma_avalon_master_readdata),                             //                                       .readdata
		.pc_dma_avalon_master_readdatavalid           (pc_dma_avalon_master_readdatavalid),                        //                                       .readdatavalid
		.pc_dma_avalon_master_write                   (pc_dma_avalon_master_write),                                //                                       .write
		.pc_dma_avalon_master_writedata               (pc_dma_avalon_master_writedata),                            //                                       .writedata
		.driver_sd_avalon_slave_0_address             (mm_interconnect_0_driver_sd_avalon_slave_0_address),        //               driver_sd_avalon_slave_0.address
		.driver_sd_avalon_slave_0_write               (mm_interconnect_0_driver_sd_avalon_slave_0_write),          //                                       .write
		.driver_sd_avalon_slave_0_read                (mm_interconnect_0_driver_sd_avalon_slave_0_read),           //                                       .read
		.driver_sd_avalon_slave_0_readdata            (mm_interconnect_0_driver_sd_avalon_slave_0_readdata),       //                                       .readdata
		.driver_sd_avalon_slave_0_writedata           (mm_interconnect_0_driver_sd_avalon_slave_0_writedata),      //                                       .writedata
		.floppy_io_address                            (mm_interconnect_0_floppy_io_address),                       //                              floppy_io.address
		.floppy_io_write                              (mm_interconnect_0_floppy_io_write),                         //                                       .write
		.floppy_io_read                               (mm_interconnect_0_floppy_io_read),                          //                                       .read
		.floppy_io_readdata                           (mm_interconnect_0_floppy_io_readdata),                      //                                       .readdata
		.floppy_io_writedata                          (mm_interconnect_0_floppy_io_writedata),                     //                                       .writedata
		.floppy_mgmt_address                          (mm_interconnect_0_floppy_mgmt_address),                     //                            floppy_mgmt.address
		.floppy_mgmt_write                            (mm_interconnect_0_floppy_mgmt_write),                       //                                       .write
		.floppy_mgmt_writedata                        (mm_interconnect_0_floppy_mgmt_writedata),                   //                                       .writedata
		.floppy_sd_slave_address                      (mm_interconnect_0_floppy_sd_slave_address),                 //                        floppy_sd_slave.address
		.floppy_sd_slave_write                        (mm_interconnect_0_floppy_sd_slave_write),                   //                                       .write
		.floppy_sd_slave_read                         (mm_interconnect_0_floppy_sd_slave_read),                    //                                       .read
		.floppy_sd_slave_readdata                     (mm_interconnect_0_floppy_sd_slave_readdata),                //                                       .readdata
		.floppy_sd_slave_writedata                    (mm_interconnect_0_floppy_sd_slave_writedata),               //                                       .writedata
		.hdd_io_address                               (mm_interconnect_0_hdd_io_address),                          //                                 hdd_io.address
		.hdd_io_write                                 (mm_interconnect_0_hdd_io_write),                            //                                       .write
		.hdd_io_read                                  (mm_interconnect_0_hdd_io_read),                             //                                       .read
		.hdd_io_readdata                              (mm_interconnect_0_hdd_io_readdata),                         //                                       .readdata
		.hdd_io_writedata                             (mm_interconnect_0_hdd_io_writedata),                        //                                       .writedata
		.hdd_io_byteenable                            (mm_interconnect_0_hdd_io_byteenable),                       //                                       .byteenable
		.hdd_mgmt_address                             (mm_interconnect_0_hdd_mgmt_address),                        //                               hdd_mgmt.address
		.hdd_mgmt_write                               (mm_interconnect_0_hdd_mgmt_write),                          //                                       .write
		.hdd_mgmt_writedata                           (mm_interconnect_0_hdd_mgmt_writedata),                      //                                       .writedata
		.hdd_sd_slave_address                         (mm_interconnect_0_hdd_sd_slave_address),                    //                           hdd_sd_slave.address
		.hdd_sd_slave_write                           (mm_interconnect_0_hdd_sd_slave_write),                      //                                       .write
		.hdd_sd_slave_read                            (mm_interconnect_0_hdd_sd_slave_read),                       //                                       .read
		.hdd_sd_slave_readdata                        (mm_interconnect_0_hdd_sd_slave_readdata),                   //                                       .readdata
		.hdd_sd_slave_writedata                       (mm_interconnect_0_hdd_sd_slave_writedata),                  //                                       .writedata
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.nios2_jtag_debug_module_address              (mm_interconnect_0_nios2_jtag_debug_module_address),         //                nios2_jtag_debug_module.address
		.nios2_jtag_debug_module_write                (mm_interconnect_0_nios2_jtag_debug_module_write),           //                                       .write
		.nios2_jtag_debug_module_read                 (mm_interconnect_0_nios2_jtag_debug_module_read),            //                                       .read
		.nios2_jtag_debug_module_readdata             (mm_interconnect_0_nios2_jtag_debug_module_readdata),        //                                       .readdata
		.nios2_jtag_debug_module_writedata            (mm_interconnect_0_nios2_jtag_debug_module_writedata),       //                                       .writedata
		.nios2_jtag_debug_module_byteenable           (mm_interconnect_0_nios2_jtag_debug_module_byteenable),      //                                       .byteenable
		.nios2_jtag_debug_module_waitrequest          (mm_interconnect_0_nios2_jtag_debug_module_waitrequest),     //                                       .waitrequest
		.nios2_jtag_debug_module_debugaccess          (mm_interconnect_0_nios2_jtag_debug_module_debugaccess),     //                                       .debugaccess
		.onchip_for_nios2_s1_address                  (mm_interconnect_0_onchip_for_nios2_s1_address),             //                    onchip_for_nios2_s1.address
		.onchip_for_nios2_s1_write                    (mm_interconnect_0_onchip_for_nios2_s1_write),               //                                       .write
		.onchip_for_nios2_s1_readdata                 (mm_interconnect_0_onchip_for_nios2_s1_readdata),            //                                       .readdata
		.onchip_for_nios2_s1_writedata                (mm_interconnect_0_onchip_for_nios2_s1_writedata),           //                                       .writedata
		.onchip_for_nios2_s1_byteenable               (mm_interconnect_0_onchip_for_nios2_s1_byteenable),          //                                       .byteenable
		.onchip_for_nios2_s1_chipselect               (mm_interconnect_0_onchip_for_nios2_s1_chipselect),          //                                       .chipselect
		.onchip_for_nios2_s1_clken                    (mm_interconnect_0_onchip_for_nios2_s1_clken),               //                                       .clken
		.pc_bus_ctrl_address                          (mm_interconnect_0_pc_bus_ctrl_address),                     //                            pc_bus_ctrl.address
		.pc_bus_ctrl_write                            (mm_interconnect_0_pc_bus_ctrl_write),                       //                                       .write
		.pc_bus_ctrl_writedata                        (mm_interconnect_0_pc_bus_ctrl_writedata),                   //                                       .writedata
		.pc_dma_master_address                        (mm_interconnect_0_pc_dma_master_address),                   //                          pc_dma_master.address
		.pc_dma_master_write                          (mm_interconnect_0_pc_dma_master_write),                     //                                       .write
		.pc_dma_master_read                           (mm_interconnect_0_pc_dma_master_read),                      //                                       .read
		.pc_dma_master_readdata                       (mm_interconnect_0_pc_dma_master_readdata),                  //                                       .readdata
		.pc_dma_master_writedata                      (mm_interconnect_0_pc_dma_master_writedata),                 //                                       .writedata
		.pc_dma_page_address                          (mm_interconnect_0_pc_dma_page_address),                     //                            pc_dma_page.address
		.pc_dma_page_write                            (mm_interconnect_0_pc_dma_page_write),                       //                                       .write
		.pc_dma_page_read                             (mm_interconnect_0_pc_dma_page_read),                        //                                       .read
		.pc_dma_page_readdata                         (mm_interconnect_0_pc_dma_page_readdata),                    //                                       .readdata
		.pc_dma_page_writedata                        (mm_interconnect_0_pc_dma_page_writedata),                   //                                       .writedata
		.pc_dma_slave_address                         (mm_interconnect_0_pc_dma_slave_address),                    //                           pc_dma_slave.address
		.pc_dma_slave_write                           (mm_interconnect_0_pc_dma_slave_write),                      //                                       .write
		.pc_dma_slave_read                            (mm_interconnect_0_pc_dma_slave_read),                       //                                       .read
		.pc_dma_slave_readdata                        (mm_interconnect_0_pc_dma_slave_readdata),                   //                                       .readdata
		.pc_dma_slave_writedata                       (mm_interconnect_0_pc_dma_slave_writedata),                  //                                       .writedata
		.pic_master_address                           (mm_interconnect_0_pic_master_address),                      //                             pic_master.address
		.pic_master_write                             (mm_interconnect_0_pic_master_write),                        //                                       .write
		.pic_master_read                              (mm_interconnect_0_pic_master_read),                         //                                       .read
		.pic_master_readdata                          (mm_interconnect_0_pic_master_readdata),                     //                                       .readdata
		.pic_master_writedata                         (mm_interconnect_0_pic_master_writedata),                    //                                       .writedata
		.pic_slave_address                            (mm_interconnect_0_pic_slave_address),                       //                              pic_slave.address
		.pic_slave_write                              (mm_interconnect_0_pic_slave_write),                         //                                       .write
		.pic_slave_read                               (mm_interconnect_0_pic_slave_read),                          //                                       .read
		.pic_slave_readdata                           (mm_interconnect_0_pic_slave_readdata),                      //                                       .readdata
		.pic_slave_writedata                          (mm_interconnect_0_pic_slave_writedata),                     //                                       .writedata
		.pio_input_s1_address                         (mm_interconnect_0_pio_input_s1_address),                    //                           pio_input_s1.address
		.pio_input_s1_write                           (mm_interconnect_0_pio_input_s1_write),                      //                                       .write
		.pio_input_s1_readdata                        (mm_interconnect_0_pio_input_s1_readdata),                   //                                       .readdata
		.pio_input_s1_writedata                       (mm_interconnect_0_pio_input_s1_writedata),                  //                                       .writedata
		.pio_input_s1_chipselect                      (mm_interconnect_0_pio_input_s1_chipselect),                 //                                       .chipselect
		.pio_output_s1_address                        (mm_interconnect_0_pio_output_s1_address),                   //                          pio_output_s1.address
		.pio_output_s1_write                          (mm_interconnect_0_pio_output_s1_write),                     //                                       .write
		.pio_output_s1_readdata                       (mm_interconnect_0_pio_output_s1_readdata),                  //                                       .readdata
		.pio_output_s1_writedata                      (mm_interconnect_0_pio_output_s1_writedata),                 //                                       .writedata
		.pio_output_s1_chipselect                     (mm_interconnect_0_pio_output_s1_chipselect),                //                                       .chipselect
		.pit_io_address                               (mm_interconnect_0_pit_io_address),                          //                                 pit_io.address
		.pit_io_write                                 (mm_interconnect_0_pit_io_write),                            //                                       .write
		.pit_io_read                                  (mm_interconnect_0_pit_io_read),                             //                                       .read
		.pit_io_readdata                              (mm_interconnect_0_pit_io_readdata),                         //                                       .readdata
		.pit_io_writedata                             (mm_interconnect_0_pit_io_writedata),                        //                                       .writedata
		.pit_mgmt_address                             (mm_interconnect_0_pit_mgmt_address),                        //                               pit_mgmt.address
		.pit_mgmt_write                               (mm_interconnect_0_pit_mgmt_write),                          //                                       .write
		.pit_mgmt_writedata                           (mm_interconnect_0_pit_mgmt_writedata),                      //                                       .writedata
		.ps2_io_address                               (mm_interconnect_0_ps2_io_address),                          //                                 ps2_io.address
		.ps2_io_write                                 (mm_interconnect_0_ps2_io_write),                            //                                       .write
		.ps2_io_read                                  (mm_interconnect_0_ps2_io_read),                             //                                       .read
		.ps2_io_readdata                              (mm_interconnect_0_ps2_io_readdata),                         //                                       .readdata
		.ps2_io_writedata                             (mm_interconnect_0_ps2_io_writedata),                        //                                       .writedata
		.ps2_sysctl_address                           (mm_interconnect_0_ps2_sysctl_address),                      //                             ps2_sysctl.address
		.ps2_sysctl_write                             (mm_interconnect_0_ps2_sysctl_write),                        //                                       .write
		.ps2_sysctl_read                              (mm_interconnect_0_ps2_sysctl_read),                         //                                       .read
		.ps2_sysctl_readdata                          (mm_interconnect_0_ps2_sysctl_readdata),                     //                                       .readdata
		.ps2_sysctl_writedata                         (mm_interconnect_0_ps2_sysctl_writedata),                    //                                       .writedata
		.rtc_io_address                               (mm_interconnect_0_rtc_io_address),                          //                                 rtc_io.address
		.rtc_io_write                                 (mm_interconnect_0_rtc_io_write),                            //                                       .write
		.rtc_io_read                                  (mm_interconnect_0_rtc_io_read),                             //                                       .read
		.rtc_io_readdata                              (mm_interconnect_0_rtc_io_readdata),                         //                                       .readdata
		.rtc_io_writedata                             (mm_interconnect_0_rtc_io_writedata),                        //                                       .writedata
		.rtc_mgmt_address                             (mm_interconnect_0_rtc_mgmt_address),                        //                               rtc_mgmt.address
		.rtc_mgmt_write                               (mm_interconnect_0_rtc_mgmt_write),                          //                                       .write
		.rtc_mgmt_writedata                           (mm_interconnect_0_rtc_mgmt_writedata),                      //                                       .writedata
		.sdram_s1_address                             (mm_interconnect_0_sdram_s1_address),                        //                               sdram_s1.address
		.sdram_s1_write                               (mm_interconnect_0_sdram_s1_write),                          //                                       .write
		.sdram_s1_read                                (mm_interconnect_0_sdram_s1_read),                           //                                       .read
		.sdram_s1_readdata                            (mm_interconnect_0_sdram_s1_readdata),                       //                                       .readdata
		.sdram_s1_writedata                           (mm_interconnect_0_sdram_s1_writedata),                      //                                       .writedata
		.sdram_s1_byteenable                          (mm_interconnect_0_sdram_s1_byteenable),                     //                                       .byteenable
		.sdram_s1_readdatavalid                       (mm_interconnect_0_sdram_s1_readdatavalid),                  //                                       .readdatavalid
		.sdram_s1_waitrequest                         (mm_interconnect_0_sdram_s1_waitrequest),                    //                                       .waitrequest
		.sdram_s1_chipselect                          (mm_interconnect_0_sdram_s1_chipselect),                     //                                       .chipselect
		.sound_fm_address                             (mm_interconnect_0_sound_fm_address),                        //                               sound_fm.address
		.sound_fm_write                               (mm_interconnect_0_sound_fm_write),                          //                                       .write
		.sound_fm_read                                (mm_interconnect_0_sound_fm_read),                           //                                       .read
		.sound_fm_readdata                            (mm_interconnect_0_sound_fm_readdata),                       //                                       .readdata
		.sound_fm_writedata                           (mm_interconnect_0_sound_fm_writedata),                      //                                       .writedata
		.sound_io_address                             (mm_interconnect_0_sound_io_address),                        //                               sound_io.address
		.sound_io_write                               (mm_interconnect_0_sound_io_write),                          //                                       .write
		.sound_io_read                                (mm_interconnect_0_sound_io_read),                           //                                       .read
		.sound_io_readdata                            (mm_interconnect_0_sound_io_readdata),                       //                                       .readdata
		.sound_io_writedata                           (mm_interconnect_0_sound_io_writedata),                      //                                       .writedata
		.sound_mgmt_address                           (mm_interconnect_0_sound_mgmt_address),                      //                             sound_mgmt.address
		.sound_mgmt_write                             (mm_interconnect_0_sound_mgmt_write),                        //                                       .write
		.sound_mgmt_writedata                         (mm_interconnect_0_sound_mgmt_writedata),                    //                                       .writedata
		.vga_io_b_address                             (mm_interconnect_0_vga_io_b_address),                        //                               vga_io_b.address
		.vga_io_b_write                               (mm_interconnect_0_vga_io_b_write),                          //                                       .write
		.vga_io_b_read                                (mm_interconnect_0_vga_io_b_read),                           //                                       .read
		.vga_io_b_readdata                            (mm_interconnect_0_vga_io_b_readdata),                       //                                       .readdata
		.vga_io_b_writedata                           (mm_interconnect_0_vga_io_b_writedata),                      //                                       .writedata
		.vga_io_c_address                             (mm_interconnect_0_vga_io_c_address),                        //                               vga_io_c.address
		.vga_io_c_write                               (mm_interconnect_0_vga_io_c_write),                          //                                       .write
		.vga_io_c_read                                (mm_interconnect_0_vga_io_c_read),                           //                                       .read
		.vga_io_c_readdata                            (mm_interconnect_0_vga_io_c_readdata),                       //                                       .readdata
		.vga_io_c_writedata                           (mm_interconnect_0_vga_io_c_writedata),                      //                                       .writedata
		.vga_io_d_address                             (mm_interconnect_0_vga_io_d_address),                        //                               vga_io_d.address
		.vga_io_d_write                               (mm_interconnect_0_vga_io_d_write),                          //                                       .write
		.vga_io_d_read                                (mm_interconnect_0_vga_io_d_read),                           //                                       .read
		.vga_io_d_readdata                            (mm_interconnect_0_vga_io_d_readdata),                       //                                       .readdata
		.vga_io_d_writedata                           (mm_interconnect_0_vga_io_d_writedata),                      //                                       .writedata
		.vga_sys_address                              (mm_interconnect_0_vga_sys_address),                         //                                vga_sys.address
		.vga_sys_write                                (mm_interconnect_0_vga_sys_write),                           //                                       .write
		.vga_sys_read                                 (mm_interconnect_0_vga_sys_read),                            //                                       .read
		.vga_sys_readdata                             (mm_interconnect_0_vga_sys_readdata),                        //                                       .readdata
		.vga_sys_writedata                            (mm_interconnect_0_vga_sys_writedata)                        //                                       .writedata
	);

	system_mm_interconnect_1 mm_interconnect_1 (
		.clk_sys_clk_clk                               (clk_sys_clk),                            //                             clk_sys_clk.clk
		.clk_vga_clk_clk                               (clk_vga_clk),                            //                             clk_vga_clk.clk
		.pc_bus_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),         // pc_bus_reset_sink_reset_bridge_in_reset.reset
		.vga_reset_sink_reset_bridge_in_reset_reset    (rst_controller_001_reset_out_reset),     //    vga_reset_sink_reset_bridge_in_reset.reset
		.pc_bus_avalon_vga_master_address              (pc_bus_avalon_vga_master_address),       //                pc_bus_avalon_vga_master.address
		.pc_bus_avalon_vga_master_waitrequest          (pc_bus_avalon_vga_master_waitrequest),   //                                        .waitrequest
		.pc_bus_avalon_vga_master_burstcount           (pc_bus_avalon_vga_master_burstcount),    //                                        .burstcount
		.pc_bus_avalon_vga_master_byteenable           (pc_bus_avalon_vga_master_byteenable),    //                                        .byteenable
		.pc_bus_avalon_vga_master_read                 (pc_bus_avalon_vga_master_read),          //                                        .read
		.pc_bus_avalon_vga_master_readdata             (pc_bus_avalon_vga_master_readdata),      //                                        .readdata
		.pc_bus_avalon_vga_master_readdatavalid        (pc_bus_avalon_vga_master_readdatavalid), //                                        .readdatavalid
		.pc_bus_avalon_vga_master_write                (pc_bus_avalon_vga_master_write),         //                                        .write
		.pc_bus_avalon_vga_master_writedata            (pc_bus_avalon_vga_master_writedata),     //                                        .writedata
		.vga_mem_address                               (mm_interconnect_1_vga_mem_address),      //                                 vga_mem.address
		.vga_mem_write                                 (mm_interconnect_1_vga_mem_write),        //                                        .write
		.vga_mem_read                                  (mm_interconnect_1_vga_mem_read),         //                                        .read
		.vga_mem_readdata                              (mm_interconnect_1_vga_mem_readdata),     //                                        .readdata
		.vga_mem_writedata                             (mm_interconnect_1_vga_mem_writedata)     //                                        .writedata
	);

	system_mm_interconnect_2 mm_interconnect_2 (
		.clk_sys_clk_clk                               (clk_sys_clk),                                //                             clk_sys_clk.clk
		.ao486_reset_sink_reset_bridge_in_reset_reset  (reset_only_ao486_reset_out_reset),           //  ao486_reset_sink_reset_bridge_in_reset.reset
		.pc_bus_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),             // pc_bus_reset_sink_reset_bridge_in_reset.reset
		.ao486_avalon_memory_address                   (ao486_avalon_memory_address),                //                     ao486_avalon_memory.address
		.ao486_avalon_memory_waitrequest               (ao486_avalon_memory_waitrequest),            //                                        .waitrequest
		.ao486_avalon_memory_burstcount                (ao486_avalon_memory_burstcount),             //                                        .burstcount
		.ao486_avalon_memory_byteenable                (ao486_avalon_memory_byteenable),             //                                        .byteenable
		.ao486_avalon_memory_read                      (ao486_avalon_memory_read),                   //                                        .read
		.ao486_avalon_memory_readdata                  (ao486_avalon_memory_readdata),               //                                        .readdata
		.ao486_avalon_memory_readdatavalid             (ao486_avalon_memory_readdatavalid),          //                                        .readdatavalid
		.ao486_avalon_memory_write                     (ao486_avalon_memory_write),                  //                                        .write
		.ao486_avalon_memory_writedata                 (ao486_avalon_memory_writedata),              //                                        .writedata
		.pc_bus_mem_address                            (mm_interconnect_2_pc_bus_mem_address),       //                              pc_bus_mem.address
		.pc_bus_mem_write                              (mm_interconnect_2_pc_bus_mem_write),         //                                        .write
		.pc_bus_mem_read                               (mm_interconnect_2_pc_bus_mem_read),          //                                        .read
		.pc_bus_mem_readdata                           (mm_interconnect_2_pc_bus_mem_readdata),      //                                        .readdata
		.pc_bus_mem_writedata                          (mm_interconnect_2_pc_bus_mem_writedata),     //                                        .writedata
		.pc_bus_mem_burstcount                         (mm_interconnect_2_pc_bus_mem_burstcount),    //                                        .burstcount
		.pc_bus_mem_byteenable                         (mm_interconnect_2_pc_bus_mem_byteenable),    //                                        .byteenable
		.pc_bus_mem_readdatavalid                      (mm_interconnect_2_pc_bus_mem_readdatavalid), //                                        .readdatavalid
		.pc_bus_mem_waitrequest                        (mm_interconnect_2_pc_bus_mem_waitrequest)    //                                        .waitrequest
	);

	system_mm_interconnect_3 mm_interconnect_3 (
		.clk_sound_clk_clk                                    (clk_sound_clk),                                        //                                  clk_sound_clk.clk
		.clk_sys_clk_clk                                      (clk_sys_clk),                                          //                                    clk_sys_clk.clk
		.driver_sound_reset_sound_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),                   // driver_sound_reset_sound_reset_bridge_in_reset.reset
		.sound_reset_sink_reset_bridge_in_reset_reset         (rst_controller_reset_out_reset),                       //         sound_reset_sink_reset_bridge_in_reset.reset
		.sound_sound_master_address                           (sound_sound_master_address),                           //                             sound_sound_master.address
		.sound_sound_master_waitrequest                       (sound_sound_master_waitrequest),                       //                                               .waitrequest
		.sound_sound_master_write                             (sound_sound_master_write),                             //                                               .write
		.sound_sound_master_writedata                         (sound_sound_master_writedata),                         //                                               .writedata
		.driver_sound_sound_slave_write                       (mm_interconnect_3_driver_sound_sound_slave_write),     //                       driver_sound_sound_slave.write
		.driver_sound_sound_slave_writedata                   (mm_interconnect_3_driver_sound_sound_slave_writedata)  //                                               .writedata
	);

	system_irq_mapper irq_mapper (
		.clk           (clk_sys_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.sender_irq    (nios2_d_irq_irq)                 //    sender.irq
	);

	system_irq_mapper_001 irq_mapper_001 (
		.clk           (clk_sys_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_001_receiver0_irq),   // receiver0.irq
		.receiver1_irq (irq_mapper_001_receiver1_irq),   // receiver1.irq
		.receiver2_irq (irq_mapper_001_receiver2_irq),   // receiver2.irq
		.receiver3_irq (irq_mapper_001_receiver3_irq),   // receiver3.irq
		.receiver4_irq (irq_mapper_001_receiver4_irq),   // receiver4.irq
		.receiver5_irq (irq_mapper_001_receiver5_irq),   // receiver5.irq
		.receiver6_irq (irq_mapper_001_receiver6_irq),   // receiver6.irq
		.sender_irq    (pic_interrupt_receiver_irq)      //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_sys_reset_out_reset),          // reset_in0.reset
		.clk            (clk_sys_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (reset_sys_reset_out_reset),          // reset_in0.reset
		.clk            (clk_vga_clk),                        //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (reset_sys_reset_out_reset),          // reset_in0.reset
		.clk            (clk_sound_clk),                      //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
